<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>89.9834,4.78321,233.141,-65.9766</PageViewport>
<gate>
<ID>1</ID>
<type>AA_RAM_4x4</type>
<position>126.5,-24.5</position>
<input>
<ID>ADDRESS_0</ID>23 </input>
<input>
<ID>ADDRESS_1</ID>24 </input>
<input>
<ID>ADDRESS_2</ID>25 </input>
<input>
<ID>ADDRESS_3</ID>26 </input>
<input>
<ID>DATA_IN_0</ID>19 </input>
<input>
<ID>DATA_IN_1</ID>21 </input>
<input>
<ID>DATA_IN_2</ID>22 </input>
<input>
<ID>DATA_IN_3</ID>20 </input>
<output>
<ID>DATA_OUT_0</ID>19 </output>
<output>
<ID>DATA_OUT_1</ID>21 </output>
<output>
<ID>DATA_OUT_2</ID>22 </output>
<output>
<ID>DATA_OUT_3</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:0 1</lparam>
<lparam>Address:1 2</lparam>
<lparam>Address:2 3</lparam>
<lparam>Address:3 5</lparam>
<lparam>Address:5 8</lparam>
<lparam>Address:8 13</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>128.5,-16</position>
<gparam>LABEL_TEXT 0 1 2 3 5 8 13</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>BB_CLOCK</type>
<position>100.5,-36.5</position>
<output>
<ID>CLK</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 15</lparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>105.5,-36.5</position>
<input>
<ID>N_in0</ID>16 </input>
<input>
<ID>N_in1</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>126.5,-35.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>22 </input>
<input>
<ID>IN_3</ID>20 </input>
<output>
<ID>OUT_0</ID>23 </output>
<output>
<ID>OUT_1</ID>24 </output>
<output>
<ID>OUT_2</ID>25 </output>
<output>
<ID>OUT_3</ID>26 </output>
<input>
<ID>clock</ID>18 </input>
<input>
<ID>load</ID>17 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>16</ID>
<type>EE_VDD</type>
<position>136.5,-35.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>35</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>158,-57.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>63 </input>
<input>
<ID>IN_2</ID>64 </input>
<input>
<ID>IN_3</ID>65 </input>
<input>
<ID>IN_4</ID>66 </input>
<input>
<ID>IN_5</ID>67 </input>
<input>
<ID>IN_6</ID>68 </input>
<input>
<ID>IN_7</ID>69 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>36</ID>
<type>BE_ROM_8x8</type>
<position>146.5,-40.5</position>
<input>
<ID>ADDRESS_0</ID>23 </input>
<input>
<ID>ADDRESS_1</ID>24 </input>
<input>
<ID>ADDRESS_2</ID>25 </input>
<input>
<ID>ADDRESS_3</ID>26 </input>
<output>
<ID>DATA_OUT_0</ID>62 </output>
<output>
<ID>DATA_OUT_1</ID>63 </output>
<output>
<ID>DATA_OUT_2</ID>64 </output>
<output>
<ID>DATA_OUT_3</ID>65 </output>
<output>
<ID>DATA_OUT_4</ID>66 </output>
<output>
<ID>DATA_OUT_5</ID>67 </output>
<output>
<ID>DATA_OUT_6</ID>68 </output>
<output>
<ID>DATA_OUT_7</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:1 1</lparam>
<lparam>Address:2 2</lparam>
<lparam>Address:3 3</lparam>
<lparam>Address:4 4</lparam>
<lparam>Address:5 5</lparam>
<lparam>Address:6 6</lparam>
<lparam>Address:7 7</lparam>
<lparam>Address:8 8</lparam>
<lparam>Address:9 9</lparam>
<lparam>Address:10 16</lparam>
<lparam>Address:11 17</lparam>
<lparam>Address:12 18</lparam>
<lparam>Address:13 19</lparam>
<lparam>Address:14 20</lparam>
<lparam>Address:15 21</lparam></gate>
<gate>
<ID>46</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>138,-87.5</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>90 </input>
<input>
<ID>IN_2</ID>91 </input>
<input>
<ID>IN_3</ID>92 </input>
<input>
<ID>IN_4</ID>93 </input>
<input>
<ID>IN_5</ID>94 </input>
<input>
<ID>IN_6</ID>95 </input>
<input>
<ID>IN_7</ID>96 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>47</ID>
<type>BE_ROM_8x8</type>
<position>117.5,-59.5</position>
<input>
<ID>ADDRESS_0</ID>104 </input>
<input>
<ID>ADDRESS_1</ID>105 </input>
<input>
<ID>ADDRESS_2</ID>103 </input>
<input>
<ID>ADDRESS_3</ID>100 </input>
<input>
<ID>ADDRESS_4</ID>101 </input>
<input>
<ID>ADDRESS_5</ID>102 </input>
<input>
<ID>ADDRESS_6</ID>98 </input>
<input>
<ID>ADDRESS_7</ID>99 </input>
<output>
<ID>DATA_OUT_0</ID>89 </output>
<output>
<ID>DATA_OUT_1</ID>90 </output>
<output>
<ID>DATA_OUT_2</ID>91 </output>
<output>
<ID>DATA_OUT_3</ID>92 </output>
<output>
<ID>DATA_OUT_4</ID>93 </output>
<output>
<ID>DATA_OUT_5</ID>94 </output>
<output>
<ID>DATA_OUT_6</ID>95 </output>
<output>
<ID>DATA_OUT_7</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:1 1</lparam>
<lparam>Address:2 1</lparam>
<lparam>Address:3 2</lparam>
<lparam>Address:4 3</lparam>
<lparam>Address:5 5</lparam>
<lparam>Address:6 8</lparam>
<lparam>Address:7 19</lparam>
<lparam>Address:8 33</lparam>
<lparam>Address:9 52</lparam>
<lparam>Address:10 85</lparam>
<lparam>Address:11 137</lparam></gate>
<gate>
<ID>48</ID>
<type>BB_CLOCK</type>
<position>91.5,-69.5</position>
<output>
<ID>CLK</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 15</lparam></gate>
<gate>
<ID>49</ID>
<type>GA_LED</type>
<position>96.5,-69.5</position>
<input>
<ID>N_in0</ID>97 </input>
<input>
<ID>N_in1</ID>149 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AE_REGISTER8</type>
<position>104,-60</position>
<output>
<ID>OUT_0</ID>104 </output>
<output>
<ID>OUT_1</ID>105 </output>
<output>
<ID>OUT_2</ID>103 </output>
<output>
<ID>OUT_3</ID>100 </output>
<output>
<ID>OUT_4</ID>101 </output>
<output>
<ID>OUT_5</ID>102 </output>
<output>
<ID>OUT_6</ID>98 </output>
<output>
<ID>OUT_7</ID>99 </output>
<input>
<ID>clear</ID>148 </input>
<input>
<ID>clock</ID>149 </input>
<input>
<ID>count_enable</ID>109 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>55</ID>
<type>EE_VDD</type>
<position>104,-51</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_AND2</type>
<position>108,-68</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-36.5,104.5,-36.5</points>
<connection>
<GID>7</GID>
<name>CLK</name></connection>
<connection>
<GID>11</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,-36.5,136.5,-36.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>load</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,-36.5,121.5,-36.5</points>
<connection>
<GID>14</GID>
<name>clock</name></connection>
<connection>
<GID>11</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-32,128,-29.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-32,125,-29.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-32,127,-29.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-32,126,-29.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-44,118.5,-26</points>
<intersection>-44 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118.5,-44,141.5,-44</points>
<connection>
<GID>36</GID>
<name>ADDRESS_0</name></connection>
<intersection>118.5 0</intersection>
<intersection>128 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118.5,-26,121.5,-26</points>
<connection>
<GID>1</GID>
<name>ADDRESS_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128,-44,128,-39</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-43,117.5,-25</points>
<intersection>-43 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-43,141.5,-43</points>
<connection>
<GID>36</GID>
<name>ADDRESS_1</name></connection>
<intersection>117.5 0</intersection>
<intersection>127 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>117.5,-25,121.5,-25</points>
<connection>
<GID>1</GID>
<name>ADDRESS_1</name></connection>
<intersection>117.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127,-43,127,-39</points>
<connection>
<GID>14</GID>
<name>OUT_1</name></connection>
<intersection>-43 1</intersection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-42,116.5,-24</points>
<intersection>-42 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-42,141.5,-42</points>
<connection>
<GID>36</GID>
<name>ADDRESS_2</name></connection>
<intersection>116.5 0</intersection>
<intersection>126 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-24,121.5,-24</points>
<connection>
<GID>1</GID>
<name>ADDRESS_2</name></connection>
<intersection>116.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>126,-42,126,-39</points>
<connection>
<GID>14</GID>
<name>OUT_2</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-41,115.5,-23</points>
<intersection>-41 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-41,141.5,-41</points>
<connection>
<GID>36</GID>
<name>ADDRESS_3</name></connection>
<intersection>115.5 0</intersection>
<intersection>125 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115.5,-23,121.5,-23</points>
<connection>
<GID>1</GID>
<name>ADDRESS_3</name></connection>
<intersection>115.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>125,-41,125,-39</points>
<connection>
<GID>14</GID>
<name>OUT_3</name></connection>
<intersection>-41 1</intersection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-60.5,150,-47.5</points>
<connection>
<GID>36</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-60.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>150,-60.5,153,-60.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-59.5,149,-47.5</points>
<connection>
<GID>36</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149,-59.5,153,-59.5</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-58.5,148,-47.5</points>
<connection>
<GID>36</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148,-58.5,153,-58.5</points>
<connection>
<GID>35</GID>
<name>IN_2</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147,-57.5,147,-47.5</points>
<connection>
<GID>36</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-57.5,153,-57.5</points>
<connection>
<GID>35</GID>
<name>IN_3</name></connection>
<intersection>147 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,-56.5,146,-47.5</points>
<connection>
<GID>36</GID>
<name>DATA_OUT_4</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>146,-56.5,153,-56.5</points>
<connection>
<GID>35</GID>
<name>IN_4</name></connection>
<intersection>146 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-55.5,145,-47.5</points>
<connection>
<GID>36</GID>
<name>DATA_OUT_5</name></connection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-55.5,153,-55.5</points>
<connection>
<GID>35</GID>
<name>IN_5</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-54.5,144,-47.5</points>
<connection>
<GID>36</GID>
<name>DATA_OUT_6</name></connection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-54.5,153,-54.5</points>
<connection>
<GID>35</GID>
<name>IN_6</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-53.5,143,-47.5</points>
<connection>
<GID>36</GID>
<name>DATA_OUT_7</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-53.5,153,-53.5</points>
<connection>
<GID>35</GID>
<name>IN_7</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-90.5,121,-66.5</points>
<connection>
<GID>47</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-90.5,133,-90.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-89.5,120,-66.5</points>
<connection>
<GID>47</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-89.5,133,-89.5</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-88.5,119,-66.5</points>
<connection>
<GID>47</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-88.5,133,-88.5</points>
<connection>
<GID>46</GID>
<name>IN_2</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-87.5,118,-66.5</points>
<connection>
<GID>47</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-87.5,133,-87.5</points>
<connection>
<GID>46</GID>
<name>IN_3</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-86.5,117,-66.5</points>
<connection>
<GID>47</GID>
<name>DATA_OUT_4</name></connection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,-86.5,133,-86.5</points>
<connection>
<GID>46</GID>
<name>IN_4</name></connection>
<intersection>117 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-85.5,116,-66.5</points>
<connection>
<GID>47</GID>
<name>DATA_OUT_5</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,-85.5,133,-85.5</points>
<connection>
<GID>46</GID>
<name>IN_5</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-84.5,115,-66.5</points>
<connection>
<GID>47</GID>
<name>DATA_OUT_6</name></connection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-84.5,133,-84.5</points>
<connection>
<GID>46</GID>
<name>IN_6</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-83.5,114,-66.5</points>
<connection>
<GID>47</GID>
<name>DATA_OUT_7</name></connection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-83.5,133,-83.5</points>
<connection>
<GID>46</GID>
<name>IN_7</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-69.5,95.5,-69.5</points>
<connection>
<GID>48</GID>
<name>CLK</name></connection>
<connection>
<GID>49</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-57,112.5,-57</points>
<connection>
<GID>53</GID>
<name>OUT_6</name></connection>
<connection>
<GID>47</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-56,112.5,-56</points>
<connection>
<GID>53</GID>
<name>OUT_7</name></connection>
<connection>
<GID>47</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-60,112.5,-60</points>
<connection>
<GID>53</GID>
<name>OUT_3</name></connection>
<connection>
<GID>47</GID>
<name>ADDRESS_3</name></connection>
<intersection>111.5 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>111.5,-69,111.5,-60</points>
<intersection>-69 14</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>111,-69,111.5,-69</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>111.5 13</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-59,112.5,-59</points>
<connection>
<GID>53</GID>
<name>OUT_4</name></connection>
<connection>
<GID>47</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-58,112.5,-58</points>
<connection>
<GID>53</GID>
<name>OUT_5</name></connection>
<connection>
<GID>47</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-61,112.5,-61</points>
<connection>
<GID>53</GID>
<name>OUT_2</name></connection>
<connection>
<GID>47</GID>
<name>ADDRESS_2</name></connection>
<intersection>111 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>111,-67,111,-61</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-63,112.5,-63</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<connection>
<GID>47</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-62,112.5,-62</points>
<connection>
<GID>53</GID>
<name>OUT_1</name></connection>
<connection>
<GID>47</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-54,104,-52</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<connection>
<GID>53</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-68,105,-65</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<connection>
<GID>53</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-69.5,103,-65</points>
<connection>
<GID>53</GID>
<name>clock</name></connection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-69.5,103,-69.5</points>
<connection>
<GID>49</GID>
<name>N_in1</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,92.3957,827.446,-316.595</PageViewport>
<gate>
<ID>38</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>102,-58.5</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>82 </input>
<input>
<ID>IN_3</ID>81 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>39</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>90.5,-58.5</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>87 </input>
<input>
<ID>IN_2</ID>86 </input>
<input>
<ID>IN_3</ID>85 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>40</ID>
<type>BE_ROM_8x8</type>
<position>89,-35</position>
<input>
<ID>ADDRESS_0</ID>84 </input>
<input>
<ID>ADDRESS_1</ID>83 </input>
<input>
<ID>ADDRESS_2</ID>82 </input>
<input>
<ID>ADDRESS_3</ID>81 </input>
<input>
<ID>ADDRESS_4</ID>88 </input>
<input>
<ID>ADDRESS_5</ID>87 </input>
<input>
<ID>ADDRESS_6</ID>86 </input>
<input>
<ID>ADDRESS_7</ID>85 </input>
<output>
<ID>DATA_OUT_0</ID>71 </output>
<output>
<ID>DATA_OUT_1</ID>72 </output>
<output>
<ID>DATA_OUT_2</ID>73 </output>
<output>
<ID>DATA_OUT_3</ID>74 </output>
<output>
<ID>DATA_OUT_4</ID>76 </output>
<output>
<ID>DATA_OUT_5</ID>75 </output>
<output>
<ID>DATA_OUT_6</ID>77 </output>
<output>
<ID>DATA_OUT_7</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>41</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>84,-48</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>75 </input>
<input>
<ID>IN_2</ID>77 </input>
<input>
<ID>IN_3</ID>78 </input>
<output>
<ID>OUT_0</ID>88 </output>
<output>
<ID>OUT_1</ID>87 </output>
<output>
<ID>OUT_2</ID>86 </output>
<output>
<ID>OUT_3</ID>85 </output>
<input>
<ID>clock</ID>70 </input>
<input>
<ID>load</ID>80 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>42</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>95.5,-48</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT_0</ID>84 </output>
<output>
<ID>OUT_1</ID>83 </output>
<output>
<ID>OUT_2</ID>82 </output>
<output>
<ID>OUT_3</ID>81 </output>
<input>
<ID>clock</ID>70 </input>
<input>
<ID>load</ID>80 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>43</ID>
<type>BB_CLOCK</type>
<position>67,-48.5</position>
<output>
<ID>CLK</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 15</lparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>72,-48.5</position>
<input>
<ID>N_in0</ID>79 </input>
<input>
<ID>N_in1</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>EE_VDD</type>
<position>103,-47.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-53,90.5,-53</points>
<intersection>75.5 4</intersection>
<intersection>90.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>90.5,-53,90.5,-49</points>
<connection>
<GID>42</GID>
<name>clock</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>75.5,-53,75.5,-48.5</points>
<intersection>-53 1</intersection>
<intersection>-49 5</intersection>
<intersection>-48.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>75.5,-49,79,-49</points>
<connection>
<GID>41</GID>
<name>clock</name></connection>
<intersection>75.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>73,-48.5,75.5,-48.5</points>
<connection>
<GID>44</GID>
<name>N_in1</name></connection>
<intersection>75.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-43.5,92.5,-42</points>
<connection>
<GID>40</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>97,-44.5,97,-43.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-43.5,97,-43.5</points>
<intersection>92.5 0</intersection>
<intersection>97 1</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-43.5,91.5,-42</points>
<connection>
<GID>40</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>96,-44.5,96,-43.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-43.5,96,-43.5</points>
<intersection>91.5 0</intersection>
<intersection>96 1</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-44.5,95,-43.5</points>
<connection>
<GID>42</GID>
<name>IN_2</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>90.5,-43.5,90.5,-42</points>
<connection>
<GID>40</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-43.5,95,-43.5</points>
<intersection>90.5 1</intersection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-44.5,94,-43.5</points>
<connection>
<GID>42</GID>
<name>IN_3</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>89.5,-43.5,89.5,-42</points>
<connection>
<GID>40</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-43.5,94,-43.5</points>
<intersection>89.5 1</intersection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-44.5,84.5,-43.5</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>87.5,-43.5,87.5,-42</points>
<connection>
<GID>40</GID>
<name>DATA_OUT_5</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-43.5,87.5,-43.5</points>
<intersection>84.5 0</intersection>
<intersection>87.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-44.5,85.5,-43.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>88.5,-43.5,88.5,-42</points>
<connection>
<GID>40</GID>
<name>DATA_OUT_4</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>85.5,-43.5,88.5,-43.5</points>
<intersection>85.5 0</intersection>
<intersection>88.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-44.5,83.5,-43</points>
<connection>
<GID>41</GID>
<name>IN_2</name></connection>
<intersection>-43 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>86.5,-43,86.5,-42</points>
<connection>
<GID>40</GID>
<name>DATA_OUT_6</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>83.5,-43,86.5,-43</points>
<intersection>83.5 0</intersection>
<intersection>86.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-43,85.5,-42</points>
<connection>
<GID>40</GID>
<name>DATA_OUT_7</name></connection>
<intersection>-43 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>82.5,-44.5,82.5,-43</points>
<connection>
<GID>41</GID>
<name>IN_3</name></connection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-43,85.5,-43</points>
<intersection>82.5 1</intersection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-48.5,71,-48.5</points>
<connection>
<GID>43</GID>
<name>CLK</name></connection>
<connection>
<GID>44</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,-52,103,-52</points>
<intersection>90 4</intersection>
<intersection>103 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>103,-52,103,-48.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>-52 1</intersection>
<intersection>-49 7</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>90,-52,90,-49</points>
<intersection>-52 1</intersection>
<intersection>-49 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89,-49,90,-49</points>
<connection>
<GID>41</GID>
<name>load</name></connection>
<intersection>90 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>100.5,-49,103,-49</points>
<connection>
<GID>42</GID>
<name>load</name></connection>
<intersection>103 3</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-56.5,94,-35.5</points>
<connection>
<GID>42</GID>
<name>OUT_3</name></connection>
<intersection>-56.5 1</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94,-56.5,99,-56.5</points>
<connection>
<GID>38</GID>
<name>IN_3</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-35.5,94,-35.5</points>
<connection>
<GID>40</GID>
<name>ADDRESS_3</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-57.5,95,-36.5</points>
<connection>
<GID>42</GID>
<name>OUT_2</name></connection>
<intersection>-57.5 1</intersection>
<intersection>-36.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-57.5,99,-57.5</points>
<connection>
<GID>38</GID>
<name>IN_2</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>84,-36.5,95,-36.5</points>
<connection>
<GID>40</GID>
<name>ADDRESS_2</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-58.5,96,-37.5</points>
<connection>
<GID>42</GID>
<name>OUT_1</name></connection>
<intersection>-58.5 1</intersection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96,-58.5,99,-58.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-37.5,96,-37.5</points>
<connection>
<GID>40</GID>
<name>ADDRESS_1</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-59.5,97,-38.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-59.5 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97,-59.5,99,-59.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-38.5,97,-38.5</points>
<connection>
<GID>40</GID>
<name>ADDRESS_0</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-56.5,82.5,-31.5</points>
<connection>
<GID>41</GID>
<name>OUT_3</name></connection>
<intersection>-56.5 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-56.5,87.5,-56.5</points>
<connection>
<GID>39</GID>
<name>IN_3</name></connection>
<intersection>82.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-31.5,84,-31.5</points>
<connection>
<GID>40</GID>
<name>ADDRESS_7</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-57.5,83.5,-32.5</points>
<connection>
<GID>41</GID>
<name>OUT_2</name></connection>
<intersection>-57.5 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-57.5,87.5,-57.5</points>
<connection>
<GID>39</GID>
<name>IN_2</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,-32.5,84,-32.5</points>
<connection>
<GID>40</GID>
<name>ADDRESS_6</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-58.5,84.5,-33.5</points>
<connection>
<GID>41</GID>
<name>OUT_1</name></connection>
<intersection>-58.5 1</intersection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-58.5,87.5,-58.5</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-33.5,84.5,-33.5</points>
<connection>
<GID>40</GID>
<name>ADDRESS_5</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-59.5,85.5,-34.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>-59.5 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-59.5,87.5,-59.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-34.5,85.5,-34.5</points>
<connection>
<GID>40</GID>
<name>ADDRESS_4</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,92.3957,827.446,-316.595</PageViewport></page 2>
<page 3>
<PageViewport>0,92.3957,827.446,-316.595</PageViewport></page 3>
<page 4>
<PageViewport>0,92.3957,827.446,-316.595</PageViewport></page 4>
<page 5>
<PageViewport>0,92.3957,827.446,-316.595</PageViewport></page 5>
<page 6>
<PageViewport>0,92.3957,827.446,-316.595</PageViewport></page 6>
<page 7>
<PageViewport>0,92.3957,827.446,-316.595</PageViewport></page 7>
<page 8>
<PageViewport>0,92.3957,827.446,-316.595</PageViewport></page 8>
<page 9>
<PageViewport>0,92.3957,827.446,-316.595</PageViewport></page 9></circuit>