<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-76.8872,115.987,211.145,-34.1852</PageViewport>
<gate>
<ID>26</ID>
<type>CC_PULSE</type>
<position>-3.5,17</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>27</ID>
<type>CC_PULSE</type>
<position>0.5,39.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>28</ID>
<type>CC_PULSE</type>
<position>-3.5,39.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>29</ID>
<type>CC_PULSE</type>
<position>-7.5,39.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>30</ID>
<type>CC_PULSE</type>
<position>0.5,32</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>31</ID>
<type>CC_PULSE</type>
<position>-3.5,32</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>32</ID>
<type>CC_PULSE</type>
<position>-7.5,32</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>33</ID>
<type>CC_PULSE</type>
<position>0.5,24.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>34</ID>
<type>CC_PULSE</type>
<position>-3.5,24.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>35</ID>
<type>CC_PULSE</type>
<position>-7.5,24.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>-7.5,43.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>-3.5,43.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>0.5,43.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>-7.5,36</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>-3.5,36</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>41</ID>
<type>DE_TO</type>
<position>0.5,36</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>-7.5,28.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>-3.5,28.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>0.5,28.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>-3.5,21</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>77</ID>
<type>CC_PULSE</type>
<position>10,17</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>78</ID>
<type>DE_TO</type>
<position>10,21</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,41.5,-7.5,41.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,41.5,-3.5,41.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,41.5,0.5,41.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,34,-7.5,34</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,34,-3.5,34</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>0.5,34,0.5,34</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<connection>
<GID>41</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,26.5,-7.5,26.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,26.5,-3.5,26.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,26.5,0.5,26.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<connection>
<GID>44</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,19,-3.5,19</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,19,10,19</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>1.4183,33.4778,201.669,-70.9274</PageViewport>
<gate>
<ID>56</ID>
<type>AE_FULLADDER_4BIT</type>
<position>78.5,-32</position>
<input>
<ID>IN_3</ID>199 </input>
<input>
<ID>IN_B_0</ID>199 </input>
<input>
<ID>IN_B_1</ID>110 </input>
<input>
<ID>IN_B_2</ID>106 </input>
<input>
<ID>IN_B_3</ID>85 </input>
<output>
<ID>OUT_0</ID>202 </output>
<output>
<ID>OUT_1</ID>200 </output>
<output>
<ID>OUT_2</ID>201 </output>
<output>
<ID>OUT_3</ID>203 </output>
<output>
<ID>carry_out</ID>60 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>57</ID>
<type>AE_FULLADDER_4BIT</type>
<position>78.5,-48</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>106 </input>
<input>
<ID>IN_2</ID>85 </input>
<output>
<ID>OUT_0</ID>229 </output>
<output>
<ID>OUT_1</ID>207 </output>
<output>
<ID>OUT_2</ID>206 </output>
<output>
<ID>OUT_3</ID>205 </output>
<input>
<ID>carry_in</ID>60 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_FULLADDER_4BIT</type>
<position>112,-12</position>
<input>
<ID>IN_2</ID>202 </input>
<input>
<ID>IN_3</ID>200 </input>
<input>
<ID>IN_B_1</ID>202 </input>
<input>
<ID>IN_B_2</ID>200 </input>
<input>
<ID>IN_B_3</ID>201 </input>
<output>
<ID>OUT_0</ID>214 </output>
<output>
<ID>OUT_1</ID>215 </output>
<output>
<ID>OUT_2</ID>216 </output>
<output>
<ID>OUT_3</ID>217 </output>
<output>
<ID>carry_out</ID>210 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_FULLADDER_4BIT</type>
<position>112,-29</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>203 </input>
<input>
<ID>IN_2</ID>229 </input>
<input>
<ID>IN_3</ID>207 </input>
<input>
<ID>IN_B_0</ID>203 </input>
<input>
<ID>IN_B_1</ID>229 </input>
<input>
<ID>IN_B_2</ID>207 </input>
<input>
<ID>IN_B_3</ID>206 </input>
<output>
<ID>OUT_0</ID>218 </output>
<output>
<ID>OUT_1</ID>219 </output>
<output>
<ID>OUT_2</ID>220 </output>
<output>
<ID>OUT_3</ID>221 </output>
<input>
<ID>carry_in</ID>210 </input>
<output>
<ID>carry_out</ID>212 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_FULLADDER_4BIT</type>
<position>112,-45</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>205 </input>
<input>
<ID>IN_B_0</ID>205 </input>
<output>
<ID>OUT_0</ID>222 </output>
<output>
<ID>OUT_1</ID>223 </output>
<output>
<ID>OUT_2</ID>224 </output>
<output>
<ID>OUT_3</ID>225 </output>
<input>
<ID>carry_in</ID>212 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>65</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>44,-23.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>41 </input>
<input>
<ID>IN_3</ID>40 </input>
<output>
<ID>OUT_0</ID>59 </output>
<output>
<ID>OUT_1</ID>55 </output>
<output>
<ID>OUT_2</ID>54 </output>
<output>
<ID>OUT_3</ID>53 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>66</ID>
<type>DE_OR8</type>
<position>31.5,-34.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>35 </input>
<input>
<ID>IN_3</ID>34 </input>
<input>
<ID>IN_4</ID>30 </input>
<input>
<ID>IN_5</ID>31 </input>
<input>
<ID>IN_6</ID>32 </input>
<input>
<ID>IN_7</ID>33 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>67</ID>
<type>FF_GND</type>
<position>27.5,-33</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_OR2</type>
<position>31.5,-12.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_OR4</type>
<position>31.5,-26.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>31 </input>
<input>
<ID>IN_3</ID>38 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>70</ID>
<type>AE_OR4</type>
<position>31.5,-18.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>32 </input>
<input>
<ID>IN_3</ID>43 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_OR4</type>
<position>45,-11.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>37 </input>
<input>
<ID>IN_3</ID>36 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_OR2</type>
<position>51,-5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>BB_CLOCK</type>
<position>46,-46</position>
<output>
<ID>CLK</ID>61 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>52.5,-44</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_REGISTER4</type>
<position>52.5,-31.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>54 </input>
<input>
<ID>IN_3</ID>53 </input>
<output>
<ID>OUT_0</ID>199 </output>
<output>
<ID>OUT_1</ID>110 </output>
<output>
<ID>OUT_2</ID>106 </output>
<output>
<ID>OUT_3</ID>85 </output>
<input>
<ID>clear</ID>107 </input>
<input>
<ID>clock</ID>61 </input>
<input>
<ID>load</ID>58 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>89</ID>
<type>CC_PULSE</type>
<position>-4,-7</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>90</ID>
<type>CC_PULSE</type>
<position>0,15.5</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>91</ID>
<type>CC_PULSE</type>
<position>-4,15.5</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>92</ID>
<type>CC_PULSE</type>
<position>-8,15.5</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>93</ID>
<type>CC_PULSE</type>
<position>0,8</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>94</ID>
<type>CC_PULSE</type>
<position>-4,8</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>95</ID>
<type>CC_PULSE</type>
<position>-8,8</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>96</ID>
<type>CC_PULSE</type>
<position>0,0.5</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>97</ID>
<type>CC_PULSE</type>
<position>-4,0.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>98</ID>
<type>CC_PULSE</type>
<position>-8,0.5</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>99</ID>
<type>DE_TO</type>
<position>-8,19.5</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t7</lparam></gate>
<gate>
<ID>100</ID>
<type>DE_TO</type>
<position>-4,19.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t8</lparam></gate>
<gate>
<ID>101</ID>
<type>DE_TO</type>
<position>0,19.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t9</lparam></gate>
<gate>
<ID>102</ID>
<type>DE_TO</type>
<position>-8,12</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t4</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>-4,12</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t5</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>0,12</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t6</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>-8,4.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t1</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>-4,4.5</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t2</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_TO</type>
<position>0,4.5</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t3</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>-4,-3</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t0</lparam></gate>
<gate>
<ID>109</ID>
<type>CC_PULSE</type>
<position>-12,-10</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>-12,-6</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID tCE</lparam></gate>
<gate>
<ID>112</ID>
<type>AE_OR2</type>
<position>12,-6</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AE_OR2</type>
<position>12,-10</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_OR2</type>
<position>12,-14</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>102 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AE_OR2</type>
<position>12,-18</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>AE_OR2</type>
<position>12,-22</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_OR2</type>
<position>12,-26</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR2</type>
<position>12,-30</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>98 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_OR2</type>
<position>12,-34</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_OR2</type>
<position>12,-38</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_OR2</type>
<position>12,-42</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>7,-43</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t0</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>7,-37</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t1</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>7,-33</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t2</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>7,-29</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t3</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>7,-25</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t4</lparam></gate>
<gate>
<ID>129</ID>
<type>DA_FROM</type>
<position>7,-21</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t5</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>7,-17</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t6</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>7,-13</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t7</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>7,-9</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t8</lparam></gate>
<gate>
<ID>133</ID>
<type>DA_FROM</type>
<position>7,-5</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t9</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>7,-41</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>7,-39</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>7,-35</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>137</ID>
<type>DA_FROM</type>
<position>7,-31</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>138</ID>
<type>DA_FROM</type>
<position>7,-27</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>139</ID>
<type>DA_FROM</type>
<position>7,-23</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>140</ID>
<type>DA_FROM</type>
<position>7,-19</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>141</ID>
<type>DA_FROM</type>
<position>7,-15</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>7,-11</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>7,-7</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>144</ID>
<type>DA_FROM</type>
<position>54.5,-44</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID tCE</lparam></gate>
<gate>
<ID>145</ID>
<type>AE_OR2</type>
<position>53.5,-39</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>GA_LED</type>
<position>156.5,-12.5</position>
<input>
<ID>N_in0</ID>214 </input>
<input>
<ID>N_in1</ID>111 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>156.5,-15.5</position>
<input>
<ID>N_in0</ID>215 </input>
<input>
<ID>N_in1</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>156.5,-18.5</position>
<input>
<ID>N_in0</ID>216 </input>
<input>
<ID>N_in1</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>GA_LED</type>
<position>156.5,-21.5</position>
<input>
<ID>N_in0</ID>217 </input>
<input>
<ID>N_in1</ID>114 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>GA_LED</type>
<position>156.5,-26.5</position>
<input>
<ID>N_in0</ID>218 </input>
<input>
<ID>N_in1</ID>191 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>GA_LED</type>
<position>156.5,-29.5</position>
<input>
<ID>N_in0</ID>219 </input>
<input>
<ID>N_in1</ID>192 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>GA_LED</type>
<position>156.5,-32.5</position>
<input>
<ID>N_in0</ID>220 </input>
<input>
<ID>N_in1</ID>193 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>156.5,-35.5</position>
<input>
<ID>N_in0</ID>221 </input>
<input>
<ID>N_in1</ID>194 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>GA_LED</type>
<position>156.5,-39.5</position>
<input>
<ID>N_in0</ID>222 </input>
<input>
<ID>N_in1</ID>231 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>156.5,-42.5</position>
<input>
<ID>N_in0</ID>223 </input>
<input>
<ID>N_in1</ID>232 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>GA_LED</type>
<position>156.5,-45.5</position>
<input>
<ID>N_in0</ID>224 </input>
<input>
<ID>N_in1</ID>233 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>156.5,-48.5</position>
<input>
<ID>N_in0</ID>225 </input>
<input>
<ID>N_in1</ID>234 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>97.5,-55</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>207 </input>
<input>
<ID>IN_2</ID>206 </input>
<input>
<ID>IN_3</ID>205 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>254</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>100.5,-4</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>200 </input>
<input>
<ID>IN_2</ID>201 </input>
<input>
<ID>IN_3</ID>203 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_LABEL</type>
<position>162,-12</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>259</ID>
<type>AA_LABEL</type>
<position>162,-15</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>AA_LABEL</type>
<position>162,-17.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>AA_LABEL</type>
<position>162,-20.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>160,-25.5</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>263</ID>
<type>AA_LABEL</type>
<position>159.5,-28.5</position>
<gparam>LABEL_TEXT 5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>159.5,-32</position>
<gparam>LABEL_TEXT 6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>265</ID>
<type>AA_LABEL</type>
<position>159.5,-35</position>
<gparam>LABEL_TEXT 7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>266</ID>
<type>AA_LABEL</type>
<position>160,-39</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>AA_LABEL</type>
<position>160,-42</position>
<gparam>LABEL_TEXT 9</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>268</ID>
<type>AA_LABEL</type>
<position>160,-44.5</position>
<gparam>LABEL_TEXT 10</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>AA_LABEL</type>
<position>160.5,-48</position>
<gparam>LABEL_TEXT 11</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>271</ID>
<type>AA_LABEL</type>
<position>162,-7.5</position>
<gparam>LABEL_TEXT 2 do potegi</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>273</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>194,-44.5</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>114 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>274</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>184,-44.5</position>
<input>
<ID>IN_0</ID>191 </input>
<input>
<ID>IN_1</ID>192 </input>
<input>
<ID>IN_2</ID>193 </input>
<input>
<ID>IN_3</ID>194 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>275</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>173.5,-44</position>
<input>
<ID>IN_0</ID>231 </input>
<input>
<ID>IN_1</ID>232 </input>
<input>
<ID>IN_2</ID>233 </input>
<input>
<ID>IN_3</ID>234 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>15,-38,28.5,-38</points>
<connection>
<GID>66</GID>
<name>IN_4</name></connection>
<connection>
<GID>120</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-37,24,-27.5</points>
<intersection>-37 2</intersection>
<intersection>-30 4</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24,-37,28.5,-37</points>
<connection>
<GID>66</GID>
<name>IN_5</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24,-27.5,28.5,-27.5</points>
<connection>
<GID>69</GID>
<name>IN_2</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>15,-30,24,-30</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-36,24.5,-19.5</points>
<intersection>-36 2</intersection>
<intersection>-22.5 1</intersection>
<intersection>-19.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-22.5,24.5,-22.5</points>
<intersection>15 4</intersection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-36,28.5,-36</points>
<connection>
<GID>66</GID>
<name>IN_6</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24.5,-19.5,28.5,-19.5</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>24.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-22.5,15,-22</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>-22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-35,25,-15.5</points>
<intersection>-35 2</intersection>
<intersection>-23.5 3</intersection>
<intersection>-18.5 1</intersection>
<intersection>-15.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-18.5,25,-18.5</points>
<intersection>15 5</intersection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-35,28.5,-35</points>
<connection>
<GID>66</GID>
<name>IN_7</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25,-23.5,28.5,-23.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>25,-15.5,28.5,-15.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>15,-18.5,15,-14</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-34,25.5,-6</points>
<intersection>-34 2</intersection>
<intersection>-11.5 3</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-6,25.5,-6</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-34,28.5,-34</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25.5,-11.5,28.5,-11.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-33,28.5,-31</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-34.5,37,-14.5</points>
<intersection>-34.5 8</intersection>
<intersection>-24.5 4</intersection>
<intersection>-14.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37,-24.5,41,-24.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>37,-14.5,42,-14.5</points>
<connection>
<GID>72</GID>
<name>IN_3</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>35.5,-34.5,37,-34.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-26.5,36.5,-12.5</points>
<intersection>-26.5 2</intersection>
<intersection>-23.5 1</intersection>
<intersection>-12.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-23.5,41,-23.5</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-26.5,36.5,-26.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36.5,-12.5,42,-12.5</points>
<connection>
<GID>72</GID>
<name>IN_2</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-29.5,24,-28.5</points>
<intersection>-29.5 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-28.5,24,-28.5</points>
<intersection>20.5 3</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-29.5,28.5,-29.5</points>
<connection>
<GID>69</GID>
<name>IN_3</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20.5,-34,20.5,-28.5</points>
<intersection>-34 4</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>15,-34,20.5,-34</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>20.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-25.5,24,-17.5</points>
<intersection>-25.5 2</intersection>
<intersection>-20.5 1</intersection>
<intersection>-17.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-20.5,24,-20.5</points>
<intersection>15 4</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-25.5,28.5,-25.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24,-17.5,28.5,-17.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-20.5,15,-18</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-21.5,38,-12.5</points>
<intersection>-21.5 3</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-12.5,38,-12.5</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38,-21.5,41,-21.5</points>
<connection>
<GID>65</GID>
<name>IN_3</name></connection>
<intersection>38 0</intersection>
<intersection>40 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>40,-21.5,40,-8.5</points>
<intersection>-21.5 3</intersection>
<intersection>-8.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>40,-8.5,42,-8.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>40 6</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-22.5,36.5,-18.5</points>
<intersection>-22.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-22.5,41,-22.5</points>
<connection>
<GID>65</GID>
<name>IN_2</name></connection>
<intersection>36.5 0</intersection>
<intersection>39 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-18.5,36.5,-18.5</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>39,-22.5,39,-10.5</points>
<intersection>-22.5 1</intersection>
<intersection>-10.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>39,-10.5,42,-10.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>39 5</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-16.5,24.5,-13.5</points>
<intersection>-16.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-16.5,24.5,-16.5</points>
<intersection>15 3</intersection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-13.5,28.5,-13.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,-16.5,15,-10</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>-16.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-24.5,24,-21.5</points>
<intersection>-24.5 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-24.5,24,-24.5</points>
<intersection>15 3</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-21.5,28.5,-21.5</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,-26,15,-24.5</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-42,22,-6</points>
<intersection>-42 4</intersection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22,-6,48,-6</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>15,-42,22,-42</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-29.5,42.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_3</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-29.5,48.5,-29.5</points>
<connection>
<GID>76</GID>
<name>IN_3</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-30.5,43.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_2</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-30.5,48.5,-30.5</points>
<connection>
<GID>76</GID>
<name>IN_2</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-31.5,44.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_1</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-31.5,48.5,-31.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-11.5,49,-4</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-4,49,-4</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-26.5,51.5,-15.5</points>
<connection>
<GID>76</GID>
<name>load</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-15.5,56,-15.5</points>
<intersection>51.5 0</intersection>
<intersection>56 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>56,-15.5,56,-5</points>
<intersection>-15.5 1</intersection>
<intersection>-5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-5,56,-5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>56 2</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-32.5,45.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-32.5,48.5,-32.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-40,77.5,-40</points>
<connection>
<GID>56</GID>
<name>carry_out</name></connection>
<connection>
<GID>57</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-42,46,-35.5</points>
<connection>
<GID>74</GID>
<name>CLK</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-35.5,51.5,-35.5</points>
<connection>
<GID>76</GID>
<name>clock</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-8,17.5,-8,17.5</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,17.5,-4,17.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.43359e-008,17.5,2.43359e-008,17.5</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,10,-8,10</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,10,-4,10</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<connection>
<GID>103</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-2.43359e-008,10,2.43359e-008,10</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<connection>
<GID>104</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,2.5,-8,2.5</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,2.5,-4,2.5</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.43359e-008,2.5,2.43359e-008,2.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<connection>
<GID>107</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-5,-4,-5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-8,-12,-8</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-43,9,-43</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<connection>
<GID>123</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-25,72.5,-25</points>
<intersection>56.5 11</intersection>
<intersection>72.5 12</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>56.5,-29.5,56.5,-25</points>
<connection>
<GID>76</GID>
<name>OUT_3</name></connection>
<intersection>-25 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>72.5,-30,72.5,-25</points>
<intersection>-30 13</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>61,-30,74.5,-30</points>
<connection>
<GID>56</GID>
<name>IN_B_3</name></connection>
<intersection>61 14</intersection>
<intersection>72.5 12</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>61,-52,61,-30</points>
<intersection>-52 15</intersection>
<intersection>-30 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>61,-52,74.5,-52</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<intersection>61 14</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-37,9,-37</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<connection>
<GID>125</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-33,9,-33</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<connection>
<GID>126</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-29,9,-29</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-25,9,-25</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<connection>
<GID>128</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-21,9,-21</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-17,9,-17</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-13,9,-13</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<connection>
<GID>131</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-9,9,-9</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<connection>
<GID>132</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-5,9,-5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-41,9,-41</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-39,9,-39</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<connection>
<GID>135</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-35,9,-35</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<connection>
<GID>136</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-31,9,-31</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<connection>
<GID>137</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-27,9,-27</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-23,9,-23</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-19,9,-19</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-15,9,-15</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-11,9,-11</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<connection>
<GID>142</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-7,9,-7</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<connection>
<GID>143</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-30.5,57.5,-29</points>
<intersection>-30.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-29,74.5,-29</points>
<connection>
<GID>56</GID>
<name>IN_B_2</name></connection>
<intersection>57.5 0</intersection>
<intersection>68.5 13</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-30.5,57.5,-30.5</points>
<connection>
<GID>76</GID>
<name>OUT_2</name></connection>
<intersection>57.5 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>68.5,-51,68.5,-29</points>
<intersection>-51 14</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>68.5,-51,74.5,-51</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>68.5 13</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>53.5,-36,53.5,-35.5</points>
<connection>
<GID>76</GID>
<name>clear</name></connection>
<connection>
<GID>145</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>54.5,-42,54.5,-42</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<connection>
<GID>145</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>52.5,-42,52.5,-42</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<connection>
<GID>145</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-50,63,-28</points>
<intersection>-50 9</intersection>
<intersection>-31.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-31.5,63,-31.5</points>
<connection>
<GID>76</GID>
<name>OUT_1</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-28,74.5,-28</points>
<connection>
<GID>56</GID>
<name>IN_B_1</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>63,-50,74.5,-50</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-13,158,-12.5</points>
<intersection>-13 3</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-12.5,158,-12.5</points>
<connection>
<GID>147</GID>
<name>N_in1</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>158,-13,191,-13</points>
<intersection>158 0</intersection>
<intersection>191 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>191,-45.5,191,-13</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>-13 3</intersection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,-15.5,158.5,-13</points>
<intersection>-15.5 2</intersection>
<intersection>-13 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-15.5,158.5,-15.5</points>
<connection>
<GID>148</GID>
<name>N_in1</name></connection>
<intersection>158.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>158.5,-13,191,-13</points>
<intersection>158.5 0</intersection>
<intersection>191 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>191,-44.5,191,-13</points>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<intersection>-13 3</intersection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159.5,-18.5,159.5,-13</points>
<intersection>-18.5 2</intersection>
<intersection>-13 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-18.5,159.5,-18.5</points>
<connection>
<GID>149</GID>
<name>N_in1</name></connection>
<intersection>159.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>159.5,-13,191,-13</points>
<intersection>159.5 0</intersection>
<intersection>191 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>191,-43.5,191,-13</points>
<connection>
<GID>273</GID>
<name>IN_2</name></connection>
<intersection>-13 3</intersection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160.5,-21.5,160.5,-13</points>
<intersection>-21.5 2</intersection>
<intersection>-13 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-21.5,160.5,-21.5</points>
<connection>
<GID>150</GID>
<name>N_in1</name></connection>
<intersection>160.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>160.5,-13,191,-13</points>
<intersection>160.5 0</intersection>
<intersection>191 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>191,-42.5,191,-13</points>
<connection>
<GID>273</GID>
<name>IN_3</name></connection>
<intersection>-13 3</intersection></vsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-26.5,162,-26</points>
<intersection>-26.5 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-26.5,162,-26.5</points>
<connection>
<GID>151</GID>
<name>N_in1</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162,-26,164,-26</points>
<intersection>162 0</intersection>
<intersection>164 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>164,-28,164,-26</points>
<intersection>-28 4</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>164,-28,179,-28</points>
<intersection>164 3</intersection>
<intersection>179 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>179,-45.5,179,-28</points>
<intersection>-45.5 6</intersection>
<intersection>-28 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>179,-45.5,181,-45.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>179 5</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157.5,-30.5,164,-30.5</points>
<intersection>157.5 3</intersection>
<intersection>164 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>157.5,-30.5,157.5,-29.5</points>
<connection>
<GID>152</GID>
<name>N_in1</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>164,-30.5,164,-29.5</points>
<intersection>-30.5 1</intersection>
<intersection>-29.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>164,-29.5,179,-29.5</points>
<intersection>164 4</intersection>
<intersection>179 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>179,-44.5,179,-29.5</points>
<intersection>-44.5 8</intersection>
<intersection>-29.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>179,-44.5,181,-44.5</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>179 7</intersection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-32.5,162,-28</points>
<intersection>-32.5 1</intersection>
<intersection>-28 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-32.5,162,-32.5</points>
<connection>
<GID>153</GID>
<name>N_in1</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>162,-28,179.5,-28</points>
<intersection>162 0</intersection>
<intersection>179.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>179.5,-43.5,179.5,-28</points>
<intersection>-43.5 5</intersection>
<intersection>-28 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>179.5,-43.5,181,-43.5</points>
<connection>
<GID>274</GID>
<name>IN_2</name></connection>
<intersection>179.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-35.5,163,-25</points>
<intersection>-35.5 1</intersection>
<intersection>-25 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-35.5,163,-35.5</points>
<connection>
<GID>154</GID>
<name>N_in1</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>163,-25,182,-25</points>
<intersection>163 0</intersection>
<intersection>182 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>182,-42.5,182,-25</points>
<intersection>-42.5 6</intersection>
<intersection>-25 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>181,-42.5,182,-42.5</points>
<connection>
<GID>274</GID>
<name>IN_3</name></connection>
<intersection>182 5</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-32.5,64,-27</points>
<intersection>-32.5 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-27,74.5,-27</points>
<connection>
<GID>56</GID>
<name>IN_B_0</name></connection>
<intersection>64 0</intersection>
<intersection>69 9</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-32.5,64,-32.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>69,-37,69,-27</points>
<intersection>-37 10</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>69,-37,74.5,-37</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>69 9</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-31.5,87.5,-31.5</points>
<connection>
<GID>56</GID>
<name>OUT_1</name></connection>
<intersection>87.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>87.5,-31.5,87.5,-4</points>
<intersection>-31.5 1</intersection>
<intersection>-9 6</intersection>
<intersection>-4 10</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>87.5,-9,108,-9</points>
<connection>
<GID>60</GID>
<name>IN_B_2</name></connection>
<intersection>87.5 5</intersection>
<intersection>102.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>102.5,-17,102.5,-9</points>
<intersection>-17 8</intersection>
<intersection>-9 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>102.5,-17,108,-17</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<intersection>102.5 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>87.5,-4,97.5,-4</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>87.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89,-31,108,-31</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>89 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89,-32.5,89,-3</points>
<intersection>-32.5 9</intersection>
<intersection>-31 1</intersection>
<intersection>-10 4</intersection>
<intersection>-3 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>89,-10,108,-10</points>
<connection>
<GID>60</GID>
<name>IN_B_3</name></connection>
<intersection>89 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>82.5,-32.5,89,-32.5</points>
<connection>
<GID>56</GID>
<name>OUT_2</name></connection>
<intersection>89 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>89,-3,97.5,-3</points>
<connection>
<GID>254</GID>
<name>IN_2</name></connection>
<intersection>89 3</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-30.5,86,-30.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>86 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>86,-30.5,86,-5</points>
<intersection>-30.5 1</intersection>
<intersection>-8 6</intersection>
<intersection>-5 10</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>86,-8,108,-8</points>
<connection>
<GID>60</GID>
<name>IN_B_1</name></connection>
<intersection>86 5</intersection>
<intersection>99.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>99.5,-16,99.5,-8</points>
<intersection>-16 8</intersection>
<intersection>-8 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>99.5,-16,108,-16</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>99.5 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>86,-5,97.5,-5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>86 5</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-33.5,89.5,-33.5</points>
<connection>
<GID>56</GID>
<name>OUT_3</name></connection>
<intersection>89.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>89.5,-33.5,89.5,-2</points>
<intersection>-33.5 1</intersection>
<intersection>-32 7</intersection>
<intersection>-24 5</intersection>
<intersection>-2 9</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>89.5,-24,108,-24</points>
<connection>
<GID>61</GID>
<name>IN_B_0</name></connection>
<intersection>89.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89.5,-32,108,-32</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>89.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>89.5,-2,97.5,-2</points>
<connection>
<GID>254</GID>
<name>IN_3</name></connection>
<intersection>89.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-49.5,101,-49.5</points>
<connection>
<GID>57</GID>
<name>OUT_3</name></connection>
<intersection>94.5 12</intersection>
<intersection>101 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>101,-49.5,101,-40</points>
<intersection>-49.5 1</intersection>
<intersection>-48 11</intersection>
<intersection>-40 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>101,-40,108,-40</points>
<connection>
<GID>62</GID>
<name>IN_B_0</name></connection>
<intersection>101 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>101,-48,108,-48</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>101 8</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>94.5,-53,94.5,-49.5</points>
<connection>
<GID>251</GID>
<name>IN_3</name></connection>
<intersection>-49.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-48.5,100.5,-48.5</points>
<connection>
<GID>57</GID>
<name>OUT_2</name></connection>
<intersection>92.5 12</intersection>
<intersection>100.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>100.5,-48.5,100.5,-27</points>
<intersection>-48.5 1</intersection>
<intersection>-47 11</intersection>
<intersection>-27 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>100.5,-27,108,-27</points>
<connection>
<GID>61</GID>
<name>IN_B_3</name></connection>
<intersection>100.5 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>100.5,-47,108,-47</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>100.5 8</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>92.5,-54,92.5,-48.5</points>
<intersection>-54 13</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>92.5,-54,94.5,-54</points>
<connection>
<GID>251</GID>
<name>IN_2</name></connection>
<intersection>92.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-47.5,100,-47.5</points>
<connection>
<GID>57</GID>
<name>OUT_1</name></connection>
<intersection>87.5 31</intersection>
<intersection>100 25</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>100,-47.5,100,-26</points>
<intersection>-47.5 1</intersection>
<intersection>-34 30</intersection>
<intersection>-26 26</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>100,-26,108,-26</points>
<connection>
<GID>61</GID>
<name>IN_B_2</name></connection>
<intersection>100 25</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>100,-34,108,-34</points>
<connection>
<GID>61</GID>
<name>IN_3</name></connection>
<intersection>100 25</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>87.5,-55,87.5,-47.5</points>
<intersection>-55 32</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>87.5,-55,94.5,-55</points>
<connection>
<GID>251</GID>
<name>IN_1</name></connection>
<intersection>87.5 31</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-21,111,-20</points>
<connection>
<GID>61</GID>
<name>carry_in</name></connection>
<connection>
<GID>60</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-37,111,-37</points>
<connection>
<GID>61</GID>
<name>carry_out</name></connection>
<connection>
<GID>62</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-12.5,135.5,-10.5</points>
<intersection>-12.5 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-12.5,155.5,-12.5</points>
<connection>
<GID>147</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-10.5,135.5,-10.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-15.5,135.5,-11.5</points>
<intersection>-15.5 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-15.5,155.5,-15.5</points>
<connection>
<GID>148</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-11.5,135.5,-11.5</points>
<connection>
<GID>60</GID>
<name>OUT_1</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-18.5,135.5,-12.5</points>
<intersection>-18.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-18.5,155.5,-18.5</points>
<connection>
<GID>149</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-12.5,135.5,-12.5</points>
<connection>
<GID>60</GID>
<name>OUT_2</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-21.5,135.5,-13.5</points>
<intersection>-21.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-21.5,155.5,-21.5</points>
<connection>
<GID>150</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-13.5,135.5,-13.5</points>
<connection>
<GID>60</GID>
<name>OUT_3</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-27.5,135.5,-26.5</points>
<intersection>-27.5 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-26.5,155.5,-26.5</points>
<connection>
<GID>151</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-27.5,135.5,-27.5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-29.5,135.5,-28.5</points>
<intersection>-29.5 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-29.5,155.5,-29.5</points>
<connection>
<GID>152</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-28.5,135.5,-28.5</points>
<connection>
<GID>61</GID>
<name>OUT_1</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-32.5,135.5,-29.5</points>
<intersection>-32.5 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-32.5,155.5,-32.5</points>
<connection>
<GID>153</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-29.5,135.5,-29.5</points>
<connection>
<GID>61</GID>
<name>OUT_2</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-35.5,155.5,-35.5</points>
<connection>
<GID>154</GID>
<name>N_in0</name></connection>
<intersection>116 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116,-35.5,116,-30.5</points>
<connection>
<GID>61</GID>
<name>OUT_3</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-43.5,135.5,-39.5</points>
<intersection>-43.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-39.5,155.5,-39.5</points>
<connection>
<GID>155</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-43.5,135.5,-43.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-44.5,135.5,-42.5</points>
<intersection>-44.5 2</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-42.5,155.5,-42.5</points>
<connection>
<GID>156</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-44.5,135.5,-44.5</points>
<connection>
<GID>62</GID>
<name>OUT_1</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-45.5,155.5,-45.5</points>
<connection>
<GID>157</GID>
<name>N_in0</name></connection>
<connection>
<GID>62</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-48.5,135.5,-46.5</points>
<intersection>-48.5 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-48.5,155.5,-48.5</points>
<connection>
<GID>158</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-46.5,135.5,-46.5</points>
<connection>
<GID>62</GID>
<name>OUT_3</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-46.5,95,-25</points>
<intersection>-46.5 2</intersection>
<intersection>-33 4</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-25,108,-25</points>
<connection>
<GID>61</GID>
<name>IN_B_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-46.5,95,-46.5</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>91.5 5</intersection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>95,-33,108,-33</points>
<connection>
<GID>61</GID>
<name>IN_2</name></connection>
<intersection>95 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>91.5,-56,91.5,-46.5</points>
<intersection>-56 6</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>91.5,-56,94.5,-56</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>91.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-45,167,-39.5</points>
<intersection>-45 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-39.5,167,-39.5</points>
<connection>
<GID>155</GID>
<name>N_in1</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167,-45,170.5,-45</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157.5,-44,170.5,-44</points>
<connection>
<GID>275</GID>
<name>IN_1</name></connection>
<intersection>157.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>157.5,-44,157.5,-42.5</points>
<connection>
<GID>156</GID>
<name>N_in1</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-45.5,167,-43</points>
<intersection>-45.5 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-45.5,167,-45.5</points>
<connection>
<GID>157</GID>
<name>N_in1</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167,-43,170.5,-43</points>
<connection>
<GID>275</GID>
<name>IN_2</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-48.5,167,-42</points>
<intersection>-48.5 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-48.5,167,-48.5</points>
<connection>
<GID>158</GID>
<name>N_in1</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167,-42,170.5,-42</points>
<connection>
<GID>275</GID>
<name>IN_3</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 2>
<page 3>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 3>
<page 4>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 4>
<page 5>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 5>
<page 6>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 6>
<page 7>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 7>
<page 8>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 8>
<page 9>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 9></circuit>