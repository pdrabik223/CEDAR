<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-65.2496,269.185,624.495,-90.4294</PageViewport>
<gate>
<ID>579</ID>
<type>GA_LED</type>
<position>258,82</position>
<input>
<ID>N_in0</ID>705 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>580</ID>
<type>GA_LED</type>
<position>248,82</position>
<input>
<ID>N_in0</ID>704 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>581</ID>
<type>GA_LED</type>
<position>248,95</position>
<input>
<ID>N_in0</ID>707 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>582</ID>
<type>GA_LED</type>
<position>253,75.5</position>
<input>
<ID>N_in1</ID>706 </input>
<gparam>LED_BOX -4.1,-1.1,4.1,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>583</ID>
<type>GA_LED</type>
<position>253,101.5</position>
<input>
<ID>N_in0</ID>702 </input>
<gparam>LED_BOX -4.1,-1.1,4.1,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>584</ID>
<type>DA_FROM</type>
<position>248,92</position>
<input>
<ID>IN_0</ID>707 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID 0.</lparam></gate>
<gate>
<ID>15</ID>
<type>DA_FROM</type>
<position>233,92</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>234.5,102</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID .</lparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>243,93</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>234.5,89</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID '</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>233,79</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID 2</lparam></gate>
<gate>
<ID>46</ID>
<type>DA_FROM</type>
<position>243,79</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID 3</lparam></gate>
<gate>
<ID>47</ID>
<type>DA_FROM</type>
<position>234.5,76</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ,</lparam></gate>
<gate>
<ID>57</ID>
<type>GA_LED</type>
<position>243,95.5</position>
<input>
<ID>N_in1</ID>20 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>238,89</position>
<input>
<ID>N_in1</ID>24 </input>
<gparam>LED_BOX -4.1,-1.1,4.1,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>243,82.5</position>
<input>
<ID>N_in0</ID>86 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>233,82.5</position>
<input>
<ID>N_in0</ID>85 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>65</ID>
<type>GA_LED</type>
<position>233,95.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>238,76</position>
<input>
<ID>N_in1</ID>87 </input>
<gparam>LED_BOX -4.1,-1.1,4.1,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>150</ID>
<type>GA_LED</type>
<position>238,102</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -4.1,-1.1,4.1,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>571</ID>
<type>DA_FROM</type>
<position>249.5,101.5</position>
<input>
<ID>IN_0</ID>702 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ..</lparam></gate>
<gate>
<ID>572</ID>
<type>DA_FROM</type>
<position>258,92</position>
<input>
<ID>IN_0</ID>708 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID 1.</lparam></gate>
<gate>
<ID>573</ID>
<type>DA_FROM</type>
<position>249.5,88.5</position>
<input>
<ID>IN_0</ID>703 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID '.</lparam></gate>
<gate>
<ID>574</ID>
<type>DA_FROM</type>
<position>248,78.5</position>
<input>
<ID>IN_0</ID>704 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID 2.</lparam></gate>
<gate>
<ID>575</ID>
<type>DA_FROM</type>
<position>258,78.5</position>
<input>
<ID>IN_0</ID>705 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID 3.</lparam></gate>
<gate>
<ID>576</ID>
<type>DA_FROM</type>
<position>249.5,75.5</position>
<input>
<ID>IN_0</ID>706 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ,.</lparam></gate>
<gate>
<ID>577</ID>
<type>GA_LED</type>
<position>258,95</position>
<input>
<ID>N_in0</ID>708 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>578</ID>
<type>GA_LED</type>
<position>253,88.5</position>
<input>
<ID>N_in1</ID>703 </input>
<gparam>LED_BOX -4.1,-1.1,4.1,1.1</gparam>
<gparam>angle 180</gparam></gate>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,94,233,94.5</points>
<connection>
<GID>65</GID>
<name>N_in0</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,91,243,96.5</points>
<connection>
<GID>57</GID>
<name>N_in1</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>13</ID>
<points>236.5,102,239,102</points>
<connection>
<GID>150</GID>
<name>N_in0</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>236.5,89,237,89</points>
<connection>
<GID>58</GID>
<name>N_in1</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,81,233,81.5</points>
<connection>
<GID>60</GID>
<name>N_in0</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,81,243,81.5</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>236.5,76,237,76</points>
<connection>
<GID>149</GID>
<name>N_in1</name></connection>
<connection>
<GID>47</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>702</ID>
<shape>
<hsegment>
<ID>13</ID>
<points>251.5,101.5,254,101.5</points>
<connection>
<GID>583</GID>
<name>N_in0</name></connection>
<connection>
<GID>571</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>703</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>251.5,89,252,89</points>
<intersection>251.5 5</intersection>
<intersection>252 7</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>251.5,88.5,251.5,89</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>89 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>252,88.5,252,89</points>
<connection>
<GID>578</GID>
<name>N_in1</name></connection>
<intersection>89 2</intersection></vsegment></shape></wire>
<wire>
<ID>704</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,80.5,248,81</points>
<connection>
<GID>580</GID>
<name>N_in0</name></connection>
<connection>
<GID>574</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>705</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,80.5,258,81</points>
<connection>
<GID>579</GID>
<name>N_in0</name></connection>
<connection>
<GID>575</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>706</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>251.5,75.5,252,75.5</points>
<connection>
<GID>582</GID>
<name>N_in1</name></connection>
<connection>
<GID>576</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>707</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,94,248,94</points>
<connection>
<GID>581</GID>
<name>N_in0</name></connection>
<connection>
<GID>584</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>708</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,94,258,94</points>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<connection>
<GID>577</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-12.9012,156.733,407.769,-62.5931</PageViewport>
<gate>
<ID>1</ID>
<type>AE_REGISTER8</type>
<position>128.5,-27.5</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>197 </input>
<input>
<ID>IN_2</ID>196 </input>
<input>
<ID>IN_3</ID>195 </input>
<input>
<ID>IN_4</ID>194 </input>
<input>
<ID>IN_5</ID>193 </input>
<input>
<ID>IN_6</ID>192 </input>
<input>
<ID>IN_7</ID>191 </input>
<output>
<ID>OUT_0</ID>244 </output>
<output>
<ID>OUT_1</ID>245 </output>
<output>
<ID>OUT_2</ID>246 </output>
<output>
<ID>OUT_3</ID>247 </output>
<output>
<ID>OUT_4</ID>248 </output>
<output>
<ID>OUT_5</ID>249 </output>
<output>
<ID>OUT_6</ID>250 </output>
<output>
<ID>OUT_7</ID>251 </output>
<input>
<ID>clear</ID>258 </input>
<input>
<ID>clock</ID>257 </input>
<input>
<ID>load</ID>25 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>4</ID>
<type>DA_FROM</type>
<position>118.5,-50</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>70,-23.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_SMALL_INVERTER</type>
<position>74,-23.5</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>DA_FROM</type>
<position>132,-43</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_OR2</type>
<position>137,-2.5</position>
<input>
<ID>IN_0</ID>588 </input>
<input>
<ID>IN_1</ID>586 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_SMALL_INVERTER</type>
<position>86,-23.5</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_SMALL_INVERTER</type>
<position>90,-23.5</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>78,-23.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_SMALL_INVERTER</type>
<position>82,-23.5</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>100.5,-36</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>23</ID>
<type>CC_PULSE</type>
<position>21,-21</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>25</ID>
<type>DE_TO</type>
<position>21,-17</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID -</lparam></gate>
<gate>
<ID>415</ID>
<type>AE_REGISTER8</type>
<position>139,5.5</position>
<input>
<ID>IN_0</ID>576 </input>
<input>
<ID>IN_1</ID>575 </input>
<input>
<ID>IN_2</ID>574 </input>
<input>
<ID>IN_3</ID>573 </input>
<input>
<ID>IN_4</ID>563 </input>
<input>
<ID>IN_5</ID>286 </input>
<input>
<ID>IN_6</ID>285 </input>
<input>
<ID>IN_7</ID>282 </input>
<output>
<ID>OUT_0</ID>767 </output>
<output>
<ID>OUT_1</ID>766 </output>
<output>
<ID>OUT_2</ID>765 </output>
<output>
<ID>OUT_3</ID>764 </output>
<output>
<ID>OUT_4</ID>763 </output>
<output>
<ID>OUT_5</ID>762 </output>
<output>
<ID>OUT_6</ID>761 </output>
<output>
<ID>OUT_7</ID>760 </output>
<input>
<ID>clear</ID>586 </input>
<input>
<ID>clock</ID>2 </input>
<input>
<ID>load</ID>588 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_OR4</type>
<position>121.5,-45</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>28 </input>
<input>
<ID>IN_2</ID>33 </input>
<input>
<ID>IN_3</ID>29 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>416</ID>
<type>DA_FROM</type>
<position>146,-5.5</position>
<input>
<ID>IN_0</ID>587 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>418</ID>
<type>DE_TO</type>
<position>93,-50</position>
<input>
<ID>IN_0</ID>565 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>419</ID>
<type>DE_TO</type>
<position>95,-59.5</position>
<input>
<ID>IN_0</ID>566 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SUB</lparam></gate>
<gate>
<ID>420</ID>
<type>DE_TO</type>
<position>100,-50</position>
<input>
<ID>IN_0</ID>567 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID MUL</lparam></gate>
<gate>
<ID>421</ID>
<type>DE_TO</type>
<position>103.5,-50</position>
<input>
<ID>IN_0</ID>568 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID DIV</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>122.5,-50</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID *</lparam></gate>
<gate>
<ID>423</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>169,9</position>
<input>
<ID>ENABLE_0</ID>591 </input>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>225 </input>
<input>
<ID>IN_2</ID>226 </input>
<input>
<ID>IN_3</ID>228 </input>
<input>
<ID>IN_4</ID>238 </input>
<input>
<ID>IN_5</ID>237 </input>
<input>
<ID>IN_6</ID>236 </input>
<input>
<ID>IN_7</ID>235 </input>
<output>
<ID>OUT_0</ID>584 </output>
<output>
<ID>OUT_1</ID>583 </output>
<output>
<ID>OUT_2</ID>582 </output>
<output>
<ID>OUT_3</ID>577 </output>
<output>
<ID>OUT_4</ID>580 </output>
<output>
<ID>OUT_5</ID>579 </output>
<output>
<ID>OUT_6</ID>578 </output>
<output>
<ID>OUT_7</ID>577 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>124.5,-50</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID \</lparam></gate>
<gate>
<ID>426</ID>
<type>DA_FROM</type>
<position>163,3.5</position>
<input>
<ID>IN_0</ID>591 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>120.5,-50</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID -</lparam></gate>
<gate>
<ID>428</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>153,22</position>
<input>
<ID>ENABLE_0</ID>570 </input>
<output>
<ID>OUT_0</ID>584 </output>
<output>
<ID>OUT_1</ID>583 </output>
<output>
<ID>OUT_2</ID>582 </output>
<output>
<ID>OUT_3</ID>577 </output>
<output>
<ID>OUT_4</ID>580 </output>
<output>
<ID>OUT_5</ID>579 </output>
<output>
<ID>OUT_6</ID>578 </output>
<output>
<ID>OUT_7</ID>577 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>429</ID>
<type>DE_TO</type>
<position>169.5,19</position>
<input>
<ID>IN_0</ID>570 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID MUL</lparam></gate>
<gate>
<ID>42</ID>
<type>BE_JKFF_LOW</type>
<position>86.5,-55</position>
<input>
<ID>J</ID>34 </input>
<input>
<ID>K</ID>34 </input>
<output>
<ID>Q</ID>30 </output>
<input>
<ID>clear</ID>52 </input>
<input>
<ID>clock</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>44</ID>
<type>BE_JKFF_LOW</type>
<position>86.5,-45</position>
<input>
<ID>J</ID>32 </input>
<input>
<ID>K</ID>32 </input>
<output>
<ID>Q</ID>31 </output>
<input>
<ID>clear</ID>45 </input>
<input>
<ID>clock</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>93,-53</position>
<input>
<ID>N_in0</ID>30 </input>
<input>
<ID>N_in3</ID>565 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>96.5,-53</position>
<input>
<ID>N_in2</ID>566 </input>
<input>
<ID>N_in3</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>442</ID>
<type>BM_NORX2</type>
<position>223,33.5</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>639 </input>
<output>
<ID>OUT</ID>613 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>443</ID>
<type>DE_TO</type>
<position>86,-15</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID klaw</lparam></gate>
<gate>
<ID>445</ID>
<type>AE_OR2</type>
<position>138,22.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>592 </input>
<output>
<ID>OUT</ID>588 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>446</ID>
<type>AE_OR3</type>
<position>234.5,94</position>
<input>
<ID>IN_0</ID>608 </input>
<input>
<ID>IN_1</ID>611 </input>
<input>
<ID>IN_2</ID>609 </input>
<output>
<ID>OUT</ID>607 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>447</ID>
<type>AE_SMALL_INVERTER</type>
<position>229.5,96</position>
<input>
<ID>IN_0</ID>640 </input>
<output>
<ID>OUT_0</ID>608 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>448</ID>
<type>BM_NORX2</type>
<position>228.5,93</position>
<input>
<ID>IN_0</ID>641 </input>
<input>
<ID>IN_1</ID>639 </input>
<output>
<ID>OUT</ID>611 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>449</ID>
<type>AE_SMALL_INVERTER</type>
<position>221,77</position>
<input>
<ID>IN_0</ID>640 </input>
<output>
<ID>OUT_0</ID>646 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>450</ID>
<type>AA_AND3</type>
<position>223,19</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>632 </input>
<input>
<ID>IN_2</ID>639 </input>
<output>
<ID>OUT</ID>631 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>451</ID>
<type>AE_SMALL_INVERTER</type>
<position>221,71</position>
<input>
<ID>IN_0</ID>639 </input>
<output>
<ID>OUT_0</ID>647 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>452</ID>
<type>AE_SMALL_INVERTER</type>
<position>221,67</position>
<input>
<ID>IN_0</ID>641 </input>
<output>
<ID>OUT_0</ID>648 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>453</ID>
<type>AE_OR2</type>
<position>233.5,55</position>
<input>
<ID>IN_0</ID>652 </input>
<input>
<ID>IN_1</ID>651 </input>
<output>
<ID>OUT</ID>650 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>454</ID>
<type>AA_AND2</type>
<position>227.5,52.5</position>
<input>
<ID>IN_0</ID>641 </input>
<input>
<ID>IN_1</ID>653 </input>
<output>
<ID>OUT</ID>651 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>455</ID>
<type>BM_NORX2</type>
<position>227.5,56.5</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>639 </input>
<output>
<ID>OUT</ID>652 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>456</ID>
<type>AE_SMALL_INVERTER</type>
<position>222.5,51.5</position>
<input>
<ID>IN_0</ID>639 </input>
<output>
<ID>OUT_0</ID>653 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>457</ID>
<type>AE_OR3</type>
<position>231,42.5</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>640 </input>
<input>
<ID>IN_2</ID>639 </input>
<output>
<ID>OUT</ID>654 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>94.5,-55.5</position>
<gparam>LABEL_TEXT +   -</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>458</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,44.5</position>
<input>
<ID>IN_0</ID>641 </input>
<output>
<ID>OUT_0</ID>655 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>81.5,-57</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>459</ID>
<type>AE_OR4</type>
<position>231.5,28</position>
<input>
<ID>IN_0</ID>613 </input>
<input>
<ID>IN_1</ID>629 </input>
<input>
<ID>IN_2</ID>630 </input>
<input>
<ID>IN_3</ID>631 </input>
<output>
<ID>OUT</ID>656 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>460</ID>
<type>AA_AND2</type>
<position>223,29</position>
<input>
<ID>IN_0</ID>657 </input>
<input>
<ID>IN_1</ID>641 </input>
<output>
<ID>OUT</ID>629 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>81.5,-43</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID -</lparam></gate>
<gate>
<ID>461</ID>
<type>AA_AND2</type>
<position>222.5,24.5</position>
<input>
<ID>IN_0</ID>641 </input>
<input>
<ID>IN_1</ID>658 </input>
<output>
<ID>OUT</ID>630 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>462</ID>
<type>AE_SMALL_INVERTER</type>
<position>210,30</position>
<input>
<ID>IN_0</ID>640 </input>
<output>
<ID>OUT_0</ID>657 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>463</ID>
<type>AE_SMALL_INVERTER</type>
<position>215.5,23.5</position>
<input>
<ID>IN_0</ID>639 </input>
<output>
<ID>OUT_0</ID>658 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>464</ID>
<type>AE_OR4</type>
<position>248.5,109</position>
<input>
<ID>IN_0</ID>641 </input>
<input>
<ID>IN_1</ID>636 </input>
<input>
<ID>IN_2</ID>660 </input>
<input>
<ID>IN_3</ID>661 </input>
<output>
<ID>OUT</ID>659 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>465</ID>
<type>BM_NORX2</type>
<position>242.5,108</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>639 </input>
<output>
<ID>OUT</ID>660 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>466</ID>
<type>AA_AND2</type>
<position>242.5,104</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>639 </input>
<output>
<ID>OUT</ID>661 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>467</ID>
<type>AE_SMALL_INVERTER</type>
<position>218,19</position>
<input>
<ID>IN_0</ID>641 </input>
<output>
<ID>OUT_0</ID>632 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>468</ID>
<type>AA_AND2</type>
<position>226,68</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>648 </input>
<output>
<ID>OUT</ID>645 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>469</ID>
<type>DE_TO</type>
<position>254.5,109</position>
<input>
<ID>IN_0</ID>659 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID .</lparam></gate>
<gate>
<ID>470</ID>
<type>DE_TO</type>
<position>239.5,94</position>
<input>
<ID>IN_0</ID>607 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>473</ID>
<type>DE_TO</type>
<position>239,73</position>
<input>
<ID>IN_0</ID>649 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID '</lparam></gate>
<gate>
<ID>474</ID>
<type>DE_TO</type>
<position>238.5,55</position>
<input>
<ID>IN_0</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_FULLADDER_4BIT</type>
<position>147,-20</position>
<input>
<ID>IN_0</ID>244 </input>
<input>
<ID>IN_1</ID>245 </input>
<input>
<ID>IN_2</ID>246 </input>
<input>
<ID>IN_3</ID>247 </input>
<input>
<ID>IN_B_0</ID>198 </input>
<input>
<ID>IN_B_1</ID>197 </input>
<input>
<ID>IN_B_2</ID>196 </input>
<input>
<ID>IN_B_3</ID>195 </input>
<output>
<ID>OUT_0</ID>186 </output>
<output>
<ID>OUT_1</ID>188 </output>
<output>
<ID>OUT_2</ID>187 </output>
<output>
<ID>OUT_3</ID>189 </output>
<output>
<ID>carry_out</ID>223 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>88</ID>
<type>AE_FULLADDER_4BIT</type>
<position>166.5,-17</position>
<input>
<ID>IN_1</ID>204 </input>
<input>
<ID>IN_2</ID>204 </input>
<input>
<ID>IN_B_0</ID>186 </input>
<input>
<ID>IN_B_1</ID>188 </input>
<input>
<ID>IN_B_2</ID>187 </input>
<input>
<ID>IN_B_3</ID>189 </input>
<output>
<ID>OUT_0</ID>228 </output>
<output>
<ID>OUT_1</ID>226 </output>
<output>
<ID>OUT_2</ID>225 </output>
<output>
<ID>OUT_3</ID>224 </output>
<output>
<ID>carry_out</ID>241 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>89</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>156.5,-23.5</position>
<output>
<ID>A_less_B</ID>230 </output>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_3</ID>190 </input>
<input>
<ID>IN_B_0</ID>186 </input>
<input>
<ID>IN_B_1</ID>188 </input>
<input>
<ID>IN_B_2</ID>187 </input>
<input>
<ID>IN_B_3</ID>189 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>90</ID>
<type>EE_VDD</type>
<position>151.5,-28.5</position>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>91</ID>
<type>EE_VDD</type>
<position>151.5,-25.5</position>
<output>
<ID>OUT_0</ID>199 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>481</ID>
<type>DE_TO</type>
<position>238.5,28</position>
<input>
<ID>IN_0</ID>656 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ,</lparam></gate>
<gate>
<ID>482</ID>
<type>DE_TO</type>
<position>236,42.5</position>
<input>
<ID>IN_0</ID>654 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3</lparam></gate>
<gate>
<ID>483</ID>
<type>AA_AND2</type>
<position>231,123.5</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>637 </input>
<output>
<ID>OUT</ID>635 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_FULLADDER_4BIT</type>
<position>146,-42</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>249 </input>
<input>
<ID>IN_2</ID>250 </input>
<input>
<ID>IN_3</ID>251 </input>
<input>
<ID>IN_B_0</ID>194 </input>
<input>
<ID>IN_B_1</ID>193 </input>
<input>
<ID>IN_B_2</ID>192 </input>
<input>
<ID>IN_B_3</ID>191 </input>
<output>
<ID>OUT_0</ID>211 </output>
<output>
<ID>OUT_1</ID>213 </output>
<output>
<ID>OUT_2</ID>212 </output>
<output>
<ID>OUT_3</ID>214 </output>
<input>
<ID>carry_in</ID>223 </input>
<output>
<ID>carry_out</ID>572 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>484</ID>
<type>AA_AND2</type>
<position>231,119.5</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>638 </input>
<output>
<ID>OUT</ID>634 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AE_FULLADDER_4BIT</type>
<position>185,-39</position>
<input>
<ID>IN_1</ID>222 </input>
<input>
<ID>IN_2</ID>222 </input>
<input>
<ID>IN_B_0</ID>211 </input>
<input>
<ID>IN_B_1</ID>213 </input>
<input>
<ID>IN_B_2</ID>212 </input>
<input>
<ID>IN_B_3</ID>214 </input>
<output>
<ID>OUT_0</ID>235 </output>
<output>
<ID>OUT_1</ID>236 </output>
<output>
<ID>OUT_2</ID>237 </output>
<output>
<ID>OUT_3</ID>238 </output>
<input>
<ID>carry_in</ID>241 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>96</ID>
<type>DA_FROM</type>
<position>45,-2</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>486</ID>
<type>AE_OR4</type>
<position>237.5,126.5</position>
<input>
<ID>IN_0</ID>636 </input>
<input>
<ID>IN_1</ID>642 </input>
<input>
<ID>IN_2</ID>635 </input>
<input>
<ID>IN_3</ID>634 </input>
<output>
<ID>OUT</ID>633 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>97</ID>
<type>DA_FROM</type>
<position>45,0</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>487</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>121,6</position>
<input>
<ID>ENABLE_0</ID>759 </input>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>197 </input>
<input>
<ID>IN_2</ID>196 </input>
<input>
<ID>IN_3</ID>195 </input>
<input>
<ID>IN_4</ID>194 </input>
<input>
<ID>IN_5</ID>193 </input>
<input>
<ID>IN_6</ID>192 </input>
<input>
<ID>IN_7</ID>191 </input>
<output>
<ID>OUT_0</ID>576 </output>
<output>
<ID>OUT_1</ID>575 </output>
<output>
<ID>OUT_2</ID>574 </output>
<output>
<ID>OUT_3</ID>573 </output>
<output>
<ID>OUT_4</ID>563 </output>
<output>
<ID>OUT_5</ID>286 </output>
<output>
<ID>OUT_6</ID>285 </output>
<output>
<ID>OUT_7</ID>282 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>98</ID>
<type>DA_FROM</type>
<position>45,2</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>488</ID>
<type>DA_FROM</type>
<position>121,38.5</position>
<input>
<ID>IN_0</ID>610 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>99</ID>
<type>DA_FROM</type>
<position>45,4</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>489</ID>
<type>DE_TO</type>
<position>243.5,126.5</position>
<input>
<ID>IN_0</ID>633 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>45,6</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>490</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,122.5</position>
<input>
<ID>IN_0</ID>641 </input>
<output>
<ID>OUT_0</ID>637 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>45,8</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>45,10</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>103</ID>
<type>DA_FROM</type>
<position>45,12</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>104</ID>
<type>DA_FROM</type>
<position>45,14</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>105</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>175,-45.5</position>
<output>
<ID>A_less_B</ID>571 </output>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_3</ID>54 </input>
<input>
<ID>IN_B_0</ID>211 </input>
<input>
<ID>IN_B_1</ID>213 </input>
<input>
<ID>IN_B_2</ID>212 </input>
<input>
<ID>IN_B_3</ID>214 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>106</ID>
<type>EE_VDD</type>
<position>169,-50.5</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>107</ID>
<type>AE_REGISTER8</type>
<position>79.5,-2.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>109 </input>
<input>
<ID>IN_2</ID>108 </input>
<input>
<ID>IN_3</ID>107 </input>
<output>
<ID>OUT_0</ID>175 </output>
<output>
<ID>OUT_1</ID>176 </output>
<output>
<ID>OUT_2</ID>177 </output>
<output>
<ID>OUT_3</ID>178 </output>
<input>
<ID>clock</ID>227 </input>
<input>
<ID>load</ID>227 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>108</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>220,-23</position>
<input>
<ID>IN_0</ID>228 </input>
<input>
<ID>IN_1</ID>226 </input>
<input>
<ID>IN_2</ID>225 </input>
<input>
<ID>IN_3</ID>224 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>109</ID>
<type>AE_OR2</type>
<position>161.5,-28.5</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>223 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>213,-30</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>236 </input>
<input>
<ID>IN_2</ID>237 </input>
<input>
<ID>IN_3</ID>238 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_OR2</type>
<position>180,-50.5</position>
<input>
<ID>IN_0</ID>571 </input>
<input>
<ID>IN_1</ID>572 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AI_XOR2</type>
<position>168,-47.5</position>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>EE_VDD</type>
<position>164,-48.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>115</ID>
<type>AE_OR2</type>
<position>99.5,-31</position>
<input>
<ID>IN_0</ID>256 </input>
<input>
<ID>IN_1</ID>255 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>DA_FROM</type>
<position>98.5,-36</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR2</type>
<position>127.5,-36</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>258 </input>
<output>
<ID>OUT</ID>257 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>71.5,5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>78 </input>
<input>
<ID>IN_2</ID>82 </input>
<input>
<ID>IN_3</ID>81 </input>
<output>
<ID>OUT_0</ID>110 </output>
<output>
<ID>OUT_1</ID>109 </output>
<output>
<ID>OUT_2</ID>108 </output>
<output>
<ID>OUT_3</ID>107 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>122</ID>
<type>BE_NOR4</type>
<position>79,-49</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>133 </input>
<input>
<ID>IN_2</ID>143 </input>
<input>
<ID>IN_3</ID>145 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>74,-48</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>74,-46</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>126</ID>
<type>BE_NOR4</type>
<position>75.5,-59</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>134 </input>
<input>
<ID>IN_2</ID>142 </input>
<input>
<ID>IN_3</ID>144 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>70.5,-56</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>519</ID>
<type>AE_SMALL_INVERTER</type>
<position>121,13</position>
<input>
<ID>IN_0</ID>610 </input>
<output>
<ID>OUT_0</ID>759 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>70.5,-58</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID -</lparam></gate>
<gate>
<ID>520</ID>
<type>AE_SMALL_INVERTER</type>
<position>220,118.5</position>
<input>
<ID>IN_0</ID>639 </input>
<output>
<ID>OUT_0</ID>638 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>131</ID>
<type>CC_PULSE</type>
<position>14,-13.5</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>132</ID>
<type>DE_TO</type>
<position>14,-9</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID *</lparam></gate>
<gate>
<ID>133</ID>
<type>CC_PULSE</type>
<position>14,-21</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>523</ID>
<type>BM_NORX2</type>
<position>231,127.5</position>
<input>
<ID>IN_0</ID>641 </input>
<input>
<ID>IN_1</ID>639 </input>
<output>
<ID>OUT</ID>642 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>DE_TO</type>
<position>14,-17</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID \</lparam></gate>
<gate>
<ID>524</ID>
<type>AA_AND2</type>
<position>228.5,89</position>
<input>
<ID>IN_0</ID>641 </input>
<input>
<ID>IN_1</ID>639 </input>
<output>
<ID>OUT</ID>609 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>BE_JKFF_LOW</type>
<position>87,-77.5</position>
<input>
<ID>J</ID>72 </input>
<input>
<ID>K</ID>72 </input>
<output>
<ID>Q</ID>154 </output>
<input>
<ID>clear</ID>117 </input>
<input>
<ID>clock</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>525</ID>
<type>AE_OR4</type>
<position>233,73</position>
<input>
<ID>IN_0</ID>636 </input>
<input>
<ID>IN_1</ID>643 </input>
<input>
<ID>IN_2</ID>644 </input>
<input>
<ID>IN_3</ID>645 </input>
<output>
<ID>OUT</ID>649 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>136</ID>
<type>BE_JKFF_LOW</type>
<position>87,-67.5</position>
<input>
<ID>J</ID>71 </input>
<input>
<ID>K</ID>71 </input>
<output>
<ID>Q</ID>155 </output>
<input>
<ID>clear</ID>73 </input>
<input>
<ID>clock</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>526</ID>
<type>AA_AND2</type>
<position>226,76</position>
<input>
<ID>IN_0</ID>646 </input>
<input>
<ID>IN_1</ID>641 </input>
<output>
<ID>OUT</ID>643 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>GA_LED</type>
<position>100,-53</position>
<input>
<ID>N_in1</ID>155 </input>
<input>
<ID>N_in3</ID>567 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>527</ID>
<type>AA_AND2</type>
<position>226,72</position>
<input>
<ID>IN_0</ID>641 </input>
<input>
<ID>IN_1</ID>647 </input>
<output>
<ID>OUT</ID>644 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_OR8</type>
<position>60.5,-6</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>69 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>68 </input>
<input>
<ID>IN_4</ID>64 </input>
<input>
<ID>IN_5</ID>65 </input>
<input>
<ID>IN_6</ID>66 </input>
<input>
<ID>IN_7</ID>67 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>528</ID>
<type>BM_NORX2</type>
<position>321,37.5</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>677 </input>
<output>
<ID>OUT</ID>666 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>GA_LED</type>
<position>103.5,-53</position>
<input>
<ID>N_in1</ID>154 </input>
<input>
<ID>N_in3</ID>568 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>529</ID>
<type>AE_OR3</type>
<position>333,96</position>
<input>
<ID>IN_0</ID>663 </input>
<input>
<ID>IN_1</ID>665 </input>
<input>
<ID>IN_2</ID>664 </input>
<output>
<ID>OUT</ID>662 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>140</ID>
<type>FF_GND</type>
<position>56.5,-4.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>530</ID>
<type>AE_SMALL_INVERTER</type>
<position>328,98</position>
<input>
<ID>IN_0</ID>678 </input>
<output>
<ID>OUT_0</ID>663 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>101.5,-55.5</position>
<gparam>LABEL_TEXT *   \</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>531</ID>
<type>BM_NORX2</type>
<position>327,95</position>
<input>
<ID>IN_0</ID>679 </input>
<input>
<ID>IN_1</ID>677 </input>
<output>
<ID>OUT</ID>665 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>82,-79.5</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID \</lparam></gate>
<gate>
<ID>532</ID>
<type>AE_SMALL_INVERTER</type>
<position>319.5,79</position>
<input>
<ID>IN_0</ID>678 </input>
<output>
<ID>OUT_0</ID>684 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>82,-65.5</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID *</lparam></gate>
<gate>
<ID>533</ID>
<type>AA_AND3</type>
<position>321.5,21</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>670 </input>
<input>
<ID>IN_2</ID>677 </input>
<output>
<ID>OUT</ID>669 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>144</ID>
<type>BE_NOR4</type>
<position>76.5,-71.5</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>135 </input>
<input>
<ID>IN_2</ID>138 </input>
<input>
<ID>IN_3</ID>141 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>534</ID>
<type>AE_SMALL_INVERTER</type>
<position>319.5,73</position>
<input>
<ID>IN_0</ID>677 </input>
<output>
<ID>OUT_0</ID>685 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>145</ID>
<type>AE_OR2</type>
<position>60.5,16</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>535</ID>
<type>AE_SMALL_INVERTER</type>
<position>319.5,69</position>
<input>
<ID>IN_0</ID>679 </input>
<output>
<ID>OUT_0</ID>686 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>146</ID>
<type>DA_FROM</type>
<position>71.5,-70.5</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>536</ID>
<type>AE_OR2</type>
<position>332,57</position>
<input>
<ID>IN_0</ID>690 </input>
<input>
<ID>IN_1</ID>689 </input>
<output>
<ID>OUT</ID>688 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_OR4</type>
<position>59.5,2</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>80 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>79 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>537</ID>
<type>AA_AND2</type>
<position>326,54.5</position>
<input>
<ID>IN_0</ID>679 </input>
<input>
<ID>IN_1</ID>691 </input>
<output>
<ID>OUT</ID>689 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>AE_OR4</type>
<position>59.5,10</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>80 </input>
<input>
<ID>IN_2</ID>66 </input>
<input>
<ID>IN_3</ID>84 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>538</ID>
<type>BM_NORX2</type>
<position>326,58.5</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>677 </input>
<output>
<ID>OUT</ID>690 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>539</ID>
<type>AE_SMALL_INVERTER</type>
<position>321,53.5</position>
<input>
<ID>IN_0</ID>677 </input>
<output>
<ID>OUT_0</ID>691 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>540</ID>
<type>AE_OR3</type>
<position>329.5,44.5</position>
<input>
<ID>IN_0</ID>693 </input>
<input>
<ID>IN_1</ID>678 </input>
<input>
<ID>IN_2</ID>677 </input>
<output>
<ID>OUT</ID>692 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>541</ID>
<type>AE_SMALL_INVERTER</type>
<position>324.5,46.5</position>
<input>
<ID>IN_0</ID>679 </input>
<output>
<ID>OUT_0</ID>693 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>542</ID>
<type>AE_OR4</type>
<position>330,30</position>
<input>
<ID>IN_0</ID>666 </input>
<input>
<ID>IN_1</ID>667 </input>
<input>
<ID>IN_2</ID>668 </input>
<input>
<ID>IN_3</ID>669 </input>
<output>
<ID>OUT</ID>694 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>543</ID>
<type>AA_AND2</type>
<position>321.5,31</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>679 </input>
<output>
<ID>OUT</ID>667 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>155</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>110,29</position>
<input>
<ID>IN_0</ID>92 </input>
<output>
<ID>OUT_0</ID>94 </output>
<output>
<ID>carry_out</ID>93 </output>
<input>
<ID>clear</ID>93 </input>
<input>
<ID>clock</ID>232 </input>
<input>
<ID>load</ID>5 </input>
<input>
<ID>shift_enable</ID>92 </input>
<input>
<ID>shift_left</ID>92 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>544</ID>
<type>AA_AND2</type>
<position>321,26.5</position>
<input>
<ID>IN_0</ID>679 </input>
<input>
<ID>IN_1</ID>696 </input>
<output>
<ID>OUT</ID>668 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>EE_VDD</type>
<position>109.5,33.5</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>545</ID>
<type>AE_SMALL_INVERTER</type>
<position>308.5,32</position>
<input>
<ID>IN_0</ID>678 </input>
<output>
<ID>OUT_0</ID>695 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>546</ID>
<type>AE_SMALL_INVERTER</type>
<position>314,25.5</position>
<input>
<ID>IN_0</ID>677 </input>
<output>
<ID>OUT_0</ID>696 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>547</ID>
<type>AE_OR4</type>
<position>347,111</position>
<input>
<ID>IN_0</ID>679 </input>
<input>
<ID>IN_1</ID>674 </input>
<input>
<ID>IN_2</ID>698 </input>
<input>
<ID>IN_3</ID>699 </input>
<output>
<ID>OUT</ID>697 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>159</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>128.5,12.5</position>
<input>
<ID>ENABLE_0</ID>610 </input>
<input>
<ID>IN_0</ID>577 </input>
<input>
<ID>IN_1</ID>578 </input>
<input>
<ID>IN_2</ID>579 </input>
<input>
<ID>IN_3</ID>580 </input>
<input>
<ID>IN_4</ID>577 </input>
<input>
<ID>IN_5</ID>582 </input>
<input>
<ID>IN_6</ID>583 </input>
<input>
<ID>IN_7</ID>584 </input>
<output>
<ID>OUT_0</ID>282 </output>
<output>
<ID>OUT_1</ID>285 </output>
<output>
<ID>OUT_2</ID>286 </output>
<output>
<ID>OUT_3</ID>563 </output>
<output>
<ID>OUT_4</ID>573 </output>
<output>
<ID>OUT_5</ID>574 </output>
<output>
<ID>OUT_6</ID>575 </output>
<output>
<ID>OUT_7</ID>576 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>548</ID>
<type>BM_NORX2</type>
<position>341,110</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>677 </input>
<output>
<ID>OUT</ID>698 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>AE_OR2</type>
<position>141,-2.5</position>
<input>
<ID>IN_0</ID>589 </input>
<input>
<ID>IN_1</ID>587 </input>
<output>
<ID>OUT</ID>586 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>549</ID>
<type>AA_AND2</type>
<position>341,106</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>677 </input>
<output>
<ID>OUT</ID>699 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>DA_FROM</type>
<position>140,-8.5</position>
<input>
<ID>IN_0</ID>589 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>550</ID>
<type>AE_SMALL_INVERTER</type>
<position>316.5,21</position>
<input>
<ID>IN_0</ID>679 </input>
<output>
<ID>OUT_0</ID>670 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>162</ID>
<type>AE_SMALL_INVERTER</type>
<position>133.5,26.5</position>
<input>
<ID>IN_0</ID>593 </input>
<output>
<ID>OUT_0</ID>592 </output>
<gparam>angle 0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>551</ID>
<type>AA_AND2</type>
<position>324.5,70</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>686 </input>
<output>
<ID>OUT</ID>683 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>163</ID>
<type>AE_SMALL_INVERTER</type>
<position>129.5,26.5</position>
<input>
<ID>IN_0</ID>594 </input>
<output>
<ID>OUT_0</ID>593 </output>
<gparam>angle 0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>552</ID>
<type>DE_TO</type>
<position>353,111</position>
<input>
<ID>IN_0</ID>697 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ..</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_SMALL_INVERTER</type>
<position>125.5,26.5</position>
<input>
<ID>IN_0</ID>595 </input>
<output>
<ID>OUT_0</ID>594 </output>
<gparam>angle 0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>553</ID>
<type>DE_TO</type>
<position>338,96</position>
<input>
<ID>IN_0</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1.</lparam></gate>
<gate>
<ID>165</ID>
<type>AE_SMALL_INVERTER</type>
<position>123.5,30.5</position>
<input>
<ID>IN_0</ID>610 </input>
<output>
<ID>OUT_0</ID>595 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>554</ID>
<type>DE_TO</type>
<position>337.5,75</position>
<input>
<ID>IN_0</ID>687 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID '.</lparam></gate>
<gate>
<ID>555</ID>
<type>DE_TO</type>
<position>337,57</position>
<input>
<ID>IN_0</ID>688 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2.</lparam></gate>
<gate>
<ID>556</ID>
<type>DE_TO</type>
<position>337,30</position>
<input>
<ID>IN_0</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ,.</lparam></gate>
<gate>
<ID>557</ID>
<type>DE_TO</type>
<position>334.5,44.5</position>
<input>
<ID>IN_0</ID>692 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3.</lparam></gate>
<gate>
<ID>558</ID>
<type>AA_AND2</type>
<position>329.5,125.5</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>673 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>DA_FROM</type>
<position>71.5,-68.5</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>559</ID>
<type>AA_AND2</type>
<position>329.5,121.5</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>676 </input>
<output>
<ID>OUT</ID>672 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>BE_NOR4</type>
<position>77,-82</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>136 </input>
<input>
<ID>IN_2</ID>139 </input>
<input>
<ID>IN_3</ID>140 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>561</ID>
<type>AE_OR4</type>
<position>336,128.5</position>
<input>
<ID>IN_0</ID>674 </input>
<input>
<ID>IN_1</ID>680 </input>
<input>
<ID>IN_2</ID>673 </input>
<input>
<ID>IN_3</ID>672 </input>
<output>
<ID>OUT</ID>671 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>72,-79</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>562</ID>
<type>DE_TO</type>
<position>342,128.5</position>
<input>
<ID>IN_0</ID>671 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0.</lparam></gate>
<gate>
<ID>563</ID>
<type>AE_SMALL_INVERTER</type>
<position>324.5,124.5</position>
<input>
<ID>IN_0</ID>679 </input>
<output>
<ID>OUT_0</ID>675 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>564</ID>
<type>AE_SMALL_INVERTER</type>
<position>318.5,120.5</position>
<input>
<ID>IN_0</ID>677 </input>
<output>
<ID>OUT_0</ID>676 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>72,-81</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>565</ID>
<type>BM_NORX2</type>
<position>329.5,129.5</position>
<input>
<ID>IN_0</ID>679 </input>
<input>
<ID>IN_1</ID>677 </input>
<output>
<ID>OUT</ID>680 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>566</ID>
<type>AA_AND2</type>
<position>327,91</position>
<input>
<ID>IN_0</ID>679 </input>
<input>
<ID>IN_1</ID>677 </input>
<output>
<ID>OUT</ID>664 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>71.5,-72.5</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID -</lparam></gate>
<gate>
<ID>567</ID>
<type>AE_OR4</type>
<position>331.5,75</position>
<input>
<ID>IN_0</ID>674 </input>
<input>
<ID>IN_1</ID>681 </input>
<input>
<ID>IN_2</ID>682 </input>
<input>
<ID>IN_3</ID>683 </input>
<output>
<ID>OUT</ID>687 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>45,-4</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>568</ID>
<type>AA_AND2</type>
<position>324.5,78</position>
<input>
<ID>IN_0</ID>684 </input>
<input>
<ID>IN_1</ID>679 </input>
<output>
<ID>OUT</ID>681 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>DA_FROM</type>
<position>72,-83</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID -</lparam></gate>
<gate>
<ID>569</ID>
<type>AA_AND2</type>
<position>324.5,74</position>
<input>
<ID>IN_0</ID>679 </input>
<input>
<ID>IN_1</ID>685 </input>
<output>
<ID>OUT</ID>682 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>DA_FROM</type>
<position>72,-85</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID *</lparam></gate>
<gate>
<ID>181</ID>
<type>DA_FROM</type>
<position>71.5,-74.5</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID \</lparam></gate>
<gate>
<ID>182</ID>
<type>DA_FROM</type>
<position>70.5,-60</position>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID *</lparam></gate>
<gate>
<ID>183</ID>
<type>AE_OR4</type>
<position>68.5,-6</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>78 </input>
<input>
<ID>IN_3</ID>77 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>184</ID>
<type>DA_FROM</type>
<position>74,-50</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID *</lparam></gate>
<gate>
<ID>185</ID>
<type>AE_OR2</type>
<position>75.5,-9.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>186</ID>
<type>DA_FROM</type>
<position>70.5,-62</position>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID \</lparam></gate>
<gate>
<ID>187</ID>
<type>DA_FROM</type>
<position>74,-52</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID \</lparam></gate>
<gate>
<ID>194</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>99.5,-3</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>176 </input>
<input>
<ID>IN_2</ID>177 </input>
<input>
<ID>IN_3</ID>178 </input>
<output>
<ID>OUT_0</ID>198 </output>
<output>
<ID>OUT_1</ID>197 </output>
<output>
<ID>OUT_2</ID>196 </output>
<output>
<ID>OUT_3</ID>195 </output>
<output>
<ID>carry_out</ID>120 </output>
<input>
<ID>clear</ID>254 </input>
<input>
<ID>clock</ID>232 </input>
<input>
<ID>load</ID>5 </input>
<input>
<ID>shift_enable</ID>122 </input>
<input>
<ID>shift_left</ID>181 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>196</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>129.5,-9.5</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>197 </input>
<input>
<ID>IN_2</ID>196 </input>
<input>
<ID>IN_3</ID>195 </input>
<input>
<ID>IN_4</ID>194 </input>
<input>
<ID>IN_5</ID>193 </input>
<input>
<ID>IN_6</ID>192 </input>
<input>
<ID>IN_7</ID>191 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>197</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>99.5,-16</position>
<output>
<ID>OUT_0</ID>194 </output>
<output>
<ID>OUT_1</ID>193 </output>
<output>
<ID>OUT_2</ID>192 </output>
<output>
<ID>OUT_3</ID>191 </output>
<input>
<ID>carry_in</ID>120 </input>
<input>
<ID>clear</ID>254 </input>
<input>
<ID>clock</ID>232 </input>
<input>
<ID>shift_enable</ID>122 </input>
<input>
<ID>shift_left</ID>229 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>205</ID>
<type>BB_CLOCK</type>
<position>44.5,-26</position>
<output>
<ID>CLK</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>611</ID>
<type>CC_PULSE</type>
<position>89,18.5</position>
<output>
<ID>OUT_0</ID>731 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>612</ID>
<type>CC_PULSE</type>
<position>93,41</position>
<output>
<ID>OUT_0</ID>724 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>613</ID>
<type>CC_PULSE</type>
<position>89,41</position>
<output>
<ID>OUT_0</ID>723 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>614</ID>
<type>CC_PULSE</type>
<position>85,41</position>
<output>
<ID>OUT_0</ID>722 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>615</ID>
<type>CC_PULSE</type>
<position>93,33.5</position>
<output>
<ID>OUT_0</ID>727 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>616</ID>
<type>CC_PULSE</type>
<position>89,33.5</position>
<output>
<ID>OUT_0</ID>726 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>617</ID>
<type>CC_PULSE</type>
<position>85,33.5</position>
<output>
<ID>OUT_0</ID>725 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>618</ID>
<type>CC_PULSE</type>
<position>93,26</position>
<output>
<ID>OUT_0</ID>730 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>619</ID>
<type>CC_PULSE</type>
<position>89,26</position>
<output>
<ID>OUT_0</ID>729 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>620</ID>
<type>CC_PULSE</type>
<position>85,26</position>
<output>
<ID>OUT_0</ID>728 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>621</ID>
<type>DE_TO</type>
<position>85,45</position>
<input>
<ID>IN_0</ID>722 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>622</ID>
<type>DE_TO</type>
<position>89,45</position>
<input>
<ID>IN_0</ID>723 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>623</ID>
<type>DE_TO</type>
<position>93,45</position>
<input>
<ID>IN_0</ID>724 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>624</ID>
<type>DE_TO</type>
<position>85,37.5</position>
<input>
<ID>IN_0</ID>725 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>625</ID>
<type>DE_TO</type>
<position>89,37.5</position>
<input>
<ID>IN_0</ID>726 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>237</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>52.5,-19.5</position>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUT_0</ID>167 </output>
<output>
<ID>OUT_1</ID>168 </output>
<output>
<ID>OUT_2</ID>169 </output>
<output>
<ID>OUT_3</ID>170 </output>
<output>
<ID>carry_out</ID>220 </output>
<input>
<ID>clear</ID>220 </input>
<input>
<ID>clock</ID>152 </input>
<input>
<ID>load</ID>227 </input>
<input>
<ID>shift_enable</ID>160 </input>
<input>
<ID>shift_left</ID>160 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>626</ID>
<type>DE_TO</type>
<position>93,37.5</position>
<input>
<ID>IN_0</ID>727 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>627</ID>
<type>DE_TO</type>
<position>85,30</position>
<input>
<ID>IN_0</ID>728 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>239</ID>
<type>EE_VDD</type>
<position>48,-18</position>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>628</ID>
<type>DE_TO</type>
<position>89,30</position>
<input>
<ID>IN_0</ID>729 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>629</ID>
<type>DE_TO</type>
<position>93,30</position>
<input>
<ID>IN_0</ID>730 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>630</ID>
<type>DE_TO</type>
<position>89,22.5</position>
<input>
<ID>IN_0</ID>731 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>631</ID>
<type>CC_PULSE</type>
<position>99,40.5</position>
<output>
<ID>OUT_0</ID>732 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>243</ID>
<type>AE_OR4</type>
<position>61,-19.5</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>168 </input>
<input>
<ID>IN_2</ID>169 </input>
<input>
<ID>IN_3</ID>170 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>632</ID>
<type>DE_TO</type>
<position>99,44.5</position>
<input>
<ID>IN_0</ID>732 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>633</ID>
<type>CC_PULSE</type>
<position>96,40.5</position>
<output>
<ID>OUT_0</ID>733 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>634</ID>
<type>DE_TO</type>
<position>96,45</position>
<input>
<ID>IN_0</ID>733 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID =</lparam></gate>
<gate>
<ID>635</ID>
<type>CC_PULSE</type>
<position>102,40.5</position>
<output>
<ID>OUT_0</ID>734 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>247</ID>
<type>GA_LED</type>
<position>74,-20.5</position>
<input>
<ID>N_in0</ID>206 </input>
<input>
<ID>N_in1</ID>174 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>636</ID>
<type>DE_TO</type>
<position>102,44.5</position>
<input>
<ID>IN_0</ID>734 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>249</ID>
<type>DE_TO</type>
<position>77,-20.5</position>
<input>
<ID>IN_0</ID>174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cc</lparam></gate>
<gate>
<ID>638</ID>
<type>HA_JUNC_2</type>
<position>171,64.5</position>
<input>
<ID>N_in0</ID>763 </input>
<input>
<ID>N_in1</ID>639 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>255</ID>
<type>EE_VDD</type>
<position>101.5,3</position>
<output>
<ID>OUT_0</ID>181 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>256</ID>
<type>EE_VDD</type>
<position>102.5,-9</position>
<output>
<ID>OUT_0</ID>229 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_AND2</type>
<position>70,-20.5</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>218 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>654</ID>
<type>HA_JUNC_2</type>
<position>171,65.5</position>
<input>
<ID>N_in0</ID>762 </input>
<input>
<ID>N_in1</ID>641 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>655</ID>
<type>HA_JUNC_2</type>
<position>171,67</position>
<input>
<ID>N_in0</ID>761 </input>
<input>
<ID>N_in1</ID>640 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>656</ID>
<type>HA_JUNC_2</type>
<position>171,68.5</position>
<input>
<ID>N_in0</ID>760 </input>
<input>
<ID>N_in1</ID>636 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>AE_SMALL_INVERTER</type>
<position>56.5,-26</position>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>270</ID>
<type>AE_SMALL_INVERTER</type>
<position>60.5,-26</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>661</ID>
<type>HA_JUNC_2</type>
<position>268.5,63.5</position>
<input>
<ID>N_in0</ID>767 </input>
<input>
<ID>N_in1</ID>677 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>662</ID>
<type>HA_JUNC_2</type>
<position>268.5,64.5</position>
<input>
<ID>N_in0</ID>766 </input>
<input>
<ID>N_in1</ID>679 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>663</ID>
<type>HA_JUNC_2</type>
<position>268.5,66</position>
<input>
<ID>N_in0</ID>765 </input>
<input>
<ID>N_in1</ID>678 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>664</ID>
<type>HA_JUNC_2</type>
<position>268.5,67.5</position>
<input>
<ID>N_in0</ID>764 </input>
<input>
<ID>N_in1</ID>674 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>278</ID>
<type>DA_FROM</type>
<position>99.5,8</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID cc</lparam></gate>
<gate>
<ID>291</ID>
<type>AE_SMALL_INVERTER</type>
<position>78,-26</position>
<input>
<ID>IN_0</ID>218 </input>
<output>
<ID>OUT_0</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>292</ID>
<type>AE_SMALL_INVERTER</type>
<position>82,-26</position>
<input>
<ID>IN_0</ID>231 </input>
<output>
<ID>OUT_0</ID>234 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>293</ID>
<type>AE_SMALL_INVERTER</type>
<position>86,-26</position>
<input>
<ID>IN_0</ID>234 </input>
<output>
<ID>OUT_0</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>294</ID>
<type>AE_SMALL_INVERTER</type>
<position>90,-26</position>
<input>
<ID>IN_0</ID>233 </input>
<output>
<ID>OUT_0</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>165,-48.5,165,-48.5</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137,0.5,138,0.5</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<connection>
<GID>415</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-26,58.5,-26</points>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection>
<connection>
<GID>270</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-23.5,72,-23.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>7</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-23.5,94,4.5</points>
<intersection>-23.5 1</intersection>
<intersection>4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-23.5,94,-23.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,4.5,100.5,4.5</points>
<intersection>94 0</intersection>
<intersection>98 6</intersection>
<intersection>100.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100.5,2,100.5,4.5</points>
<connection>
<GID>194</GID>
<name>load</name></connection>
<intersection>4.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>98,4.5,98,10.5</points>
<intersection>4.5 2</intersection>
<intersection>10.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>98,10.5,117,10.5</points>
<intersection>98 6</intersection>
<intersection>117 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>117,10.5,117,28</points>
<intersection>10.5 8</intersection>
<intersection>28 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>115,28,117,28</points>
<connection>
<GID>155</GID>
<name>load</name></connection>
<intersection>117 9</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-48,118.5,-48</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-23.5,88,-23.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<connection>
<GID>11</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-19,21,-19</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-23.5,80,-23.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>13</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-23.5,76,-23.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-23.5,84,-23.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-41,121.5,-21.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>-41 5</intersection>
<intersection>-21.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>121.5,-21.5,127.5,-21.5</points>
<connection>
<GID>1</GID>
<name>load</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>121.5,-41,126.5,-41</points>
<intersection>121.5 0</intersection>
<intersection>126.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>126.5,-41,126.5,-39</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-41 5</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-48,120.5,-48</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-48,124.5,-48</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89.5,-53,92,-53</points>
<connection>
<GID>42</GID>
<name>Q</name></connection>
<connection>
<GID>48</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-52,96.5,-43</points>
<connection>
<GID>50</GID>
<name>N_in3</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-43,96.5,-43</points>
<connection>
<GID>44</GID>
<name>Q</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-47,83.5,-43</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<connection>
<GID>44</GID>
<name>clock</name></connection>
<connection>
<GID>44</GID>
<name>K</name></connection>
<connection>
<GID>44</GID>
<name>J</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-48,122.5,-48</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>83.5,-57,83.5,-53</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<connection>
<GID>42</GID>
<name>clock</name></connection>
<connection>
<GID>42</GID>
<name>K</name></connection>
<connection>
<GID>42</GID>
<name>J</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-49,86.5,-49</points>
<connection>
<GID>44</GID>
<name>clear</name></connection>
<connection>
<GID>122</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79.5,-59,86.5,-59</points>
<connection>
<GID>42</GID>
<name>clear</name></connection>
<connection>
<GID>126</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>170,-50.5,171,-50.5</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<connection>
<GID>105</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>14,-11.5,14,-11</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<connection>
<GID>132</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-19,14,-19</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-9.5,51,-2</points>
<intersection>-9.5 2</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-2,51,-2</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-9.5,57.5,-9.5</points>
<connection>
<GID>138</GID>
<name>IN_4</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-8.5,51.5,2</points>
<intersection>-8.5 2</intersection>
<intersection>1 3</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,2,51.5,2</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-8.5,57.5,-8.5</points>
<connection>
<GID>138</GID>
<name>IN_5</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51.5,1,56.5,1</points>
<connection>
<GID>147</GID>
<name>IN_2</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-7.5,52,9</points>
<intersection>-7.5 2</intersection>
<intersection>6 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,6,52,6</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-7.5,57.5,-7.5</points>
<connection>
<GID>138</GID>
<name>IN_6</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52,9,56.5,9</points>
<connection>
<GID>148</GID>
<name>IN_2</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-6.5,52.5,13</points>
<intersection>-6.5 2</intersection>
<intersection>5 3</intersection>
<intersection>10 1</intersection>
<intersection>13 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,10,52.5,10</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-6.5,57.5,-6.5</points>
<connection>
<GID>138</GID>
<name>IN_7</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52.5,5,56.5,5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,13,56.5,13</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-5.5,53,17</points>
<intersection>-5.5 2</intersection>
<intersection>14 1</intersection>
<intersection>17 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,14,53,14</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-5.5,57.5,-5.5</points>
<connection>
<GID>138</GID>
<name>IN_3</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>53,17,57.5,17</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-4.5,57.5,-2.5</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<connection>
<GID>138</GID>
<name>IN_2</name></connection>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-69.5,84,-65.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<connection>
<GID>136</GID>
<name>clock</name></connection>
<connection>
<GID>136</GID>
<name>K</name></connection>
<connection>
<GID>136</GID>
<name>J</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>84,-79.5,84,-75.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<connection>
<GID>135</GID>
<name>clock</name></connection>
<connection>
<GID>135</GID>
<name>K</name></connection>
<connection>
<GID>135</GID>
<name>J</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80.5,-71.5,87,-71.5</points>
<connection>
<GID>136</GID>
<name>clear</name></connection>
<connection>
<GID>144</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-9,64.5,4</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>-9 6</intersection>
<intersection>4 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>64.5,4,68.5,4</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>64.5,-9,65.5,-9</points>
<connection>
<GID>183</GID>
<name>IN_3</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-7,64,5</points>
<intersection>-7 3</intersection>
<intersection>2 2</intersection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,5,68.5,5</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,2,64,2</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,-7,65.5,-7</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-1,51.5,0</points>
<intersection>-1 2</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,0,51.5,0</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-1,56.5,-1</points>
<connection>
<GID>147</GID>
<name>IN_3</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,3,51.5,11</points>
<intersection>3 2</intersection>
<intersection>8 1</intersection>
<intersection>11 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,8,51.5,8</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,3,56.5,3</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51.5,11,56.5,11</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,7,64.5,16</points>
<intersection>7 3</intersection>
<intersection>16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63.5,16,64.5,16</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64.5,7,68.5,7</points>
<connection>
<GID>119</GID>
<name>IN_3</name></connection>
<intersection>64.5 0</intersection>
<intersection>65.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>65.5,-3,65.5,7</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>7 3</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,6,64,10</points>
<intersection>6 1</intersection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,6,68.5,6</points>
<connection>
<GID>119</GID>
<name>IN_2</name></connection>
<intersection>64 0</intersection>
<intersection>65 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,10,64,10</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>64 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>65,-5,65,6</points>
<intersection>-5 6</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>65,-5,65.5,-5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>65 5</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,12,52,15</points>
<intersection>12 1</intersection>
<intersection>15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,12,52,12</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,15,57.5,15</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,4,51.5,7</points>
<intersection>4 1</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,4,51.5,4</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,7,56.5,7</points>
<connection>
<GID>148</GID>
<name>IN_3</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,27,115.5,32.5</points>
<intersection>27 2</intersection>
<intersection>29 6</intersection>
<intersection>32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110.5,32.5,115.5,32.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>110.5 7</intersection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,27,115.5,27</points>
<connection>
<GID>155</GID>
<name>shift_left</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>115,29,115.5,29</points>
<connection>
<GID>155</GID>
<name>shift_enable</name></connection>
<intersection>115.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>110.5,32.5,110.5,33.5</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<intersection>32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,29,106,30.5</points>
<intersection>29 1</intersection>
<intersection>30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,29,106,29</points>
<connection>
<GID>155</GID>
<name>clear</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105,30.5,106,30.5</points>
<connection>
<GID>155</GID>
<name>carry_out</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,25.5,129.5,30</points>
<intersection>25.5 2</intersection>
<intersection>30 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,25.5,129.5,25.5</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>129.5,30,139,30</points>
<intersection>129.5 0</intersection>
<intersection>139 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>139,25.5,139,30</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>30 3</intersection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>72.5,-8.5,72.5,-6</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<connection>
<GID>185</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-10.5,50.5,-4</points>
<intersection>-10.5 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-4,50.5,-4</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-10.5,72.5,-10.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-2.5,70,1</points>
<connection>
<GID>119</GID>
<name>OUT_3</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-2.5,75.5,-2.5</points>
<connection>
<GID>107</GID>
<name>IN_3</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-3.5,71,1</points>
<connection>
<GID>119</GID>
<name>OUT_2</name></connection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-3.5,75.5,-3.5</points>
<connection>
<GID>107</GID>
<name>IN_2</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-4.5,72,1</points>
<connection>
<GID>119</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-4.5,75.5,-4.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-5.5,73,1</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-5.5,75.5,-5.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-82,87,-81.5</points>
<connection>
<GID>135</GID>
<name>clear</name></connection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-82,87,-82</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>20</ID>
<points>98,-11,98,-8</points>
<connection>
<GID>197</GID>
<name>carry_in</name></connection>
<connection>
<GID>194</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>104.5,-10.5,104.5,6</points>
<intersection>-10.5 20</intersection>
<intersection>6 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>99.5,6,104.5,6</points>
<intersection>99.5 22</intersection>
<intersection>104.5 1</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>99.5,-10.5,104.5,-10.5</points>
<intersection>99.5 21</intersection>
<intersection>104.5 1</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>99.5,-11,99.5,-10.5</points>
<connection>
<GID>197</GID>
<name>shift_enable</name></connection>
<intersection>-10.5 20</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>99.5,2,99.5,6</points>
<connection>
<GID>194</GID>
<name>shift_enable</name></connection>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>6 18</intersection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-46,76,-46</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<connection>
<GID>124</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-56,72.5,-56</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<connection>
<GID>128</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-68.5,73.5,-68.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<connection>
<GID>169</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-79,74,-79</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<connection>
<GID>172</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-48,76,-48</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<connection>
<GID>123</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-58,72.5,-58</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<connection>
<GID>130</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-70.5,73.5,-70.5</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<connection>
<GID>146</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-81,74,-81</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<connection>
<GID>175</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-72.5,73.5,-72.5</points>
<connection>
<GID>144</GID>
<name>IN_2</name></connection>
<connection>
<GID>177</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-83,74,-83</points>
<connection>
<GID>171</GID>
<name>IN_2</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-85,74,-85</points>
<connection>
<GID>171</GID>
<name>IN_3</name></connection>
<connection>
<GID>180</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-74.5,73.5,-74.5</points>
<connection>
<GID>144</GID>
<name>IN_3</name></connection>
<connection>
<GID>181</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-60,72.5,-60</points>
<connection>
<GID>126</GID>
<name>IN_2</name></connection>
<connection>
<GID>182</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-50,76,-50</points>
<connection>
<GID>122</GID>
<name>IN_2</name></connection>
<connection>
<GID>184</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-62,72.5,-62</points>
<connection>
<GID>126</GID>
<name>IN_3</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-52,76,-52</points>
<connection>
<GID>122</GID>
<name>IN_3</name></connection>
<connection>
<GID>187</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>18</ID>
<points>53.5,-26,53.5,-24.5</points>
<connection>
<GID>237</GID>
<name>clock</name></connection>
<intersection>-26 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>48.5,-26,54.5,-26</points>
<connection>
<GID>205</GID>
<name>CLK</name></connection>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>53.5 18</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-75.5,105.5,-53</points>
<intersection>-75.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-75.5,105.5,-75.5</points>
<connection>
<GID>135</GID>
<name>Q</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-53,105.5,-53</points>
<connection>
<GID>139</GID>
<name>N_in1</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-65.5,102,-53</points>
<intersection>-65.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-65.5,102,-65.5</points>
<connection>
<GID>136</GID>
<name>Q</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101,-53,102,-53</points>
<connection>
<GID>137</GID>
<name>N_in1</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-18,49,-13.5</points>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49,-13.5,54.5,-13.5</points>
<intersection>49 0</intersection>
<intersection>52.5 14</intersection>
<intersection>54.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>54.5,-14.5,54.5,-13.5</points>
<connection>
<GID>237</GID>
<name>shift_left</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>52.5,-14.5,52.5,-13.5</points>
<connection>
<GID>237</GID>
<name>shift_enable</name></connection>
<intersection>-13.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-18,56.5,-16.5</points>
<intersection>-18 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-18,56.5,-18</points>
<connection>
<GID>237</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-16.5,58,-16.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-18.5,58,-18.5</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>56 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>56,-19,56,-18.5</points>
<connection>
<GID>237</GID>
<name>OUT_1</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-20.5,58,-20.5</points>
<connection>
<GID>243</GID>
<name>IN_2</name></connection>
<intersection>56 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>56,-20.5,56,-20</points>
<connection>
<GID>237</GID>
<name>OUT_2</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-23.5,56,-21</points>
<connection>
<GID>237</GID>
<name>OUT_3</name></connection>
<intersection>-23.5 12</intersection>
<intersection>-22.5 15</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>56,-23.5,68,-23.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>56,-22.5,58,-22.5</points>
<connection>
<GID>243</GID>
<name>IN_3</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,6.5,135,6.5</points>
<connection>
<GID>415</GID>
<name>IN_4</name></connection>
<connection>
<GID>487</GID>
<name>OUT_4</name></connection>
<intersection>128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128,6.5,128,10.5</points>
<connection>
<GID>159</GID>
<name>OUT_3</name></connection>
<intersection>6.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-20.5,75,-20.5</points>
<connection>
<GID>247</GID>
<name>N_in1</name></connection>
<connection>
<GID>249</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-5.5,91.5,-1.5</points>
<intersection>-5.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-5.5,91.5,-5.5</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-1.5,96,-1.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-52,93,-52</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<connection>
<GID>48</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-4.5,87,-2</points>
<intersection>-4.5 1</intersection>
<intersection>-2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-4.5,87,-4.5</points>
<connection>
<GID>107</GID>
<name>OUT_1</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87,-2,96,-2</points>
<intersection>87 0</intersection>
<intersection>96 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>96,-2.5,96,-2</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>-2 2</intersection></vsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-57.5,95,-54</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-54,96.5,-54</points>
<connection>
<GID>50</GID>
<name>N_in2</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-3.5,96,-3.5</points>
<connection>
<GID>194</GID>
<name>IN_2</name></connection>
<connection>
<GID>107</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-52,100,-52</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<connection>
<GID>137</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-4.5,88.5,-2.5</points>
<intersection>-4.5 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-2.5,88.5,-2.5</points>
<connection>
<GID>107</GID>
<name>OUT_3</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-4.5,96,-4.5</points>
<connection>
<GID>194</GID>
<name>IN_3</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-52,103.5,-52</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<connection>
<GID>139</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,2,101.5,2</points>
<connection>
<GID>194</GID>
<name>shift_left</name></connection>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>153,21,169.5,21</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>153 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>153,17,153,21</points>
<connection>
<GID>428</GID>
<name>ENABLE_0</name></connection>
<intersection>21 0</intersection></vsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>177,-53.5,179,-53.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<connection>
<GID>105</GID>
<name>A_less_B</name></connection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-54,145,-50</points>
<connection>
<GID>94</GID>
<name>carry_out</name></connection>
<intersection>-54 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>181,-54,181,-53.5</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>145,-54,181,-54</points>
<intersection>145 0</intersection>
<intersection>181 1</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,5.5,135,5.5</points>
<connection>
<GID>415</GID>
<name>IN_3</name></connection>
<connection>
<GID>487</GID>
<name>OUT_3</name></connection>
<intersection>129 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>129,5.5,129,10.5</points>
<connection>
<GID>159</GID>
<name>OUT_4</name></connection>
<intersection>5.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,4.5,135,4.5</points>
<connection>
<GID>415</GID>
<name>IN_2</name></connection>
<connection>
<GID>487</GID>
<name>OUT_2</name></connection>
<intersection>130 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>130,4.5,130,10.5</points>
<connection>
<GID>159</GID>
<name>OUT_5</name></connection>
<intersection>4.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,3.5,135,3.5</points>
<connection>
<GID>415</GID>
<name>IN_1</name></connection>
<connection>
<GID>487</GID>
<name>OUT_1</name></connection>
<intersection>131 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>131,3.5,131,10.5</points>
<connection>
<GID>159</GID>
<name>OUT_6</name></connection>
<intersection>3.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-18.5,152.5,-18.5</points>
<connection>
<GID>89</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<intersection>151 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>151,-18.5,151,-12</points>
<intersection>-18.5 1</intersection>
<intersection>-12 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>151,-12,162.5,-12</points>
<connection>
<GID>88</GID>
<name>IN_B_0</name></connection>
<intersection>151 6</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,2.5,135,2.5</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<connection>
<GID>487</GID>
<name>OUT_0</name></connection>
<intersection>132 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>132,2.5,132,10.5</points>
<connection>
<GID>159</GID>
<name>OUT_7</name></connection>
<intersection>2.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-20.5,152.5,-20.5</points>
<connection>
<GID>89</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>87</GID>
<name>OUT_2</name></connection>
<intersection>152 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>152,-20.5,152,-14</points>
<intersection>-20.5 1</intersection>
<intersection>-14 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>152,-14,162.5,-14</points>
<connection>
<GID>88</GID>
<name>IN_B_2</name></connection>
<intersection>152 6</intersection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,5.5,146,18.5</points>
<intersection>5.5 2</intersection>
<intersection>18 1</intersection>
<intersection>18.5 16</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,18,146,18</points>
<intersection>125 18</intersection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>146,5.5,167,5.5</points>
<connection>
<GID>423</GID>
<name>OUT_7</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>146,18.5,168,18.5</points>
<connection>
<GID>428</GID>
<name>OUT_7</name></connection>
<intersection>146 0</intersection>
<intersection>168 19</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>125,14.5,125,18</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>18 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>168,18.5,168,22.5</points>
<intersection>18.5 16</intersection>
<intersection>22.5 26</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>148,9.5,148,22.5</points>
<intersection>9.5 22</intersection>
<intersection>16 21</intersection>
<intersection>22.5 26</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>129,16,148,16</points>
<intersection>129 28</intersection>
<intersection>148 20</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>148,9.5,167,9.5</points>
<connection>
<GID>423</GID>
<name>OUT_3</name></connection>
<intersection>148 20</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>148,22.5,168,22.5</points>
<connection>
<GID>428</GID>
<name>OUT_3</name></connection>
<intersection>148 20</intersection>
<intersection>168 19</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>129,14.5,129,16</points>
<connection>
<GID>159</GID>
<name>IN_4</name></connection>
<intersection>16 21</intersection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-19.5,152.5,-19.5</points>
<connection>
<GID>89</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>87</GID>
<name>OUT_1</name></connection>
<intersection>151.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>151.5,-19.5,151.5,-13</points>
<intersection>-19.5 1</intersection>
<intersection>-13 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>151.5,-13,162.5,-13</points>
<connection>
<GID>88</GID>
<name>IN_B_1</name></connection>
<intersection>151.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,6.5,146.5,19.5</points>
<intersection>6.5 2</intersection>
<intersection>17.5 1</intersection>
<intersection>19.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,17.5,146.5,17.5</points>
<intersection>126 8</intersection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>146.5,6.5,167,6.5</points>
<connection>
<GID>423</GID>
<name>OUT_6</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>146.5,19.5,151,19.5</points>
<connection>
<GID>428</GID>
<name>OUT_6</name></connection>
<intersection>146.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>126,14.5,126,17.5</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-21.5,152.5,-21.5</points>
<connection>
<GID>89</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>87</GID>
<name>OUT_3</name></connection>
<intersection>152.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>152.5,-21.5,152.5,-15</points>
<intersection>-21.5 1</intersection>
<intersection>-15 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>152.5,-15,162.5,-15</points>
<connection>
<GID>88</GID>
<name>IN_B_3</name></connection>
<intersection>152.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,-28.5,152.5,-28.5</points>
<connection>
<GID>89</GID>
<name>IN_3</name></connection>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>579</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147,7.5,147,20.5</points>
<intersection>7.5 2</intersection>
<intersection>17 1</intersection>
<intersection>20.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,17,147,17</points>
<intersection>127 3</intersection>
<intersection>147 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147,7.5,167,7.5</points>
<connection>
<GID>423</GID>
<name>OUT_5</name></connection>
<intersection>147 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>127,14.5,127,17</points>
<connection>
<GID>159</GID>
<name>IN_2</name></connection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>147,20.5,151,20.5</points>
<connection>
<GID>428</GID>
<name>OUT_5</name></connection>
<intersection>147 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-17.5,107,-5.5</points>
<intersection>-17.5 2</intersection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-5.5,124.5,-5.5</points>
<connection>
<GID>196</GID>
<name>IN_7</name></connection>
<intersection>107 0</intersection>
<intersection>117.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-17.5,107,-17.5</points>
<connection>
<GID>197</GID>
<name>OUT_3</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>117.5,-40,117.5,9.5</points>
<intersection>-40 6</intersection>
<intersection>-23.5 4</intersection>
<intersection>-5.5 1</intersection>
<intersection>9.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>117.5,-23.5,124.5,-23.5</points>
<connection>
<GID>1</GID>
<name>IN_7</name></connection>
<intersection>117.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>117.5,-40,142,-40</points>
<connection>
<GID>94</GID>
<name>IN_B_3</name></connection>
<intersection>117.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>117.5,9.5,119,9.5</points>
<connection>
<GID>487</GID>
<name>IN_7</name></connection>
<intersection>117.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>580</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,8.5,147.5,21.5</points>
<intersection>8.5 2</intersection>
<intersection>16.5 1</intersection>
<intersection>21.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,16.5,147.5,16.5</points>
<intersection>128 3</intersection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,8.5,167,8.5</points>
<connection>
<GID>423</GID>
<name>OUT_4</name></connection>
<intersection>147.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128,14.5,128,16.5</points>
<connection>
<GID>159</GID>
<name>IN_3</name></connection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>147.5,21.5,151,21.5</points>
<connection>
<GID>428</GID>
<name>OUT_4</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-16.5,106.5,-6.5</points>
<intersection>-16.5 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-6.5,124.5,-6.5</points>
<connection>
<GID>196</GID>
<name>IN_6</name></connection>
<intersection>106.5 0</intersection>
<intersection>116.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-16.5,106.5,-16.5</points>
<connection>
<GID>197</GID>
<name>OUT_2</name></connection>
<intersection>106.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116.5,-39,116.5,8.5</points>
<intersection>-39 6</intersection>
<intersection>-24.5 4</intersection>
<intersection>-6.5 1</intersection>
<intersection>8.5 10</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>116.5,-24.5,124.5,-24.5</points>
<connection>
<GID>1</GID>
<name>IN_6</name></connection>
<intersection>116.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>116.5,-39,142,-39</points>
<connection>
<GID>94</GID>
<name>IN_B_2</name></connection>
<intersection>116.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>116.5,8.5,119,8.5</points>
<connection>
<GID>487</GID>
<name>IN_6</name></connection>
<intersection>116.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,10.5,148.5,23.5</points>
<intersection>10.5 1</intersection>
<intersection>15.5 2</intersection>
<intersection>23.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148.5,10.5,167,10.5</points>
<connection>
<GID>423</GID>
<name>OUT_2</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>130,15.5,148.5,15.5</points>
<intersection>130 8</intersection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>148.5,23.5,151,23.5</points>
<connection>
<GID>428</GID>
<name>OUT_2</name></connection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>130,14.5,130,15.5</points>
<connection>
<GID>159</GID>
<name>IN_5</name></connection>
<intersection>15.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-15.5,106,-7.5</points>
<intersection>-15.5 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-7.5,124.5,-7.5</points>
<connection>
<GID>196</GID>
<name>IN_5</name></connection>
<intersection>106 0</intersection>
<intersection>115.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-15.5,106,-15.5</points>
<connection>
<GID>197</GID>
<name>OUT_1</name></connection>
<intersection>106 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115.5,-38,115.5,7.5</points>
<intersection>-38 6</intersection>
<intersection>-25.5 4</intersection>
<intersection>-7.5 1</intersection>
<intersection>7.5 10</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>115.5,-25.5,124.5,-25.5</points>
<connection>
<GID>1</GID>
<name>IN_5</name></connection>
<intersection>115.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>115.5,-38,142,-38</points>
<connection>
<GID>94</GID>
<name>IN_B_1</name></connection>
<intersection>115.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>115.5,7.5,119,7.5</points>
<connection>
<GID>487</GID>
<name>IN_5</name></connection>
<intersection>115.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,11.5,149,24.5</points>
<intersection>11.5 1</intersection>
<intersection>15 2</intersection>
<intersection>24.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149,11.5,167,11.5</points>
<connection>
<GID>423</GID>
<name>OUT_1</name></connection>
<intersection>149 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,15,149,15</points>
<intersection>131 9</intersection>
<intersection>149 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>149,24.5,151,24.5</points>
<connection>
<GID>428</GID>
<name>OUT_1</name></connection>
<intersection>149 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>131,14.5,131,15</points>
<connection>
<GID>159</GID>
<name>IN_6</name></connection>
<intersection>15 2</intersection></vsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-14.5,105.5,-8.5</points>
<intersection>-14.5 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-8.5,124.5,-8.5</points>
<connection>
<GID>196</GID>
<name>IN_4</name></connection>
<intersection>105.5 0</intersection>
<intersection>114.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-14.5,105.5,-14.5</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114.5,-37,114.5,6.5</points>
<intersection>-37 8</intersection>
<intersection>-26.5 4</intersection>
<intersection>-8.5 1</intersection>
<intersection>6.5 12</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>114.5,-26.5,124.5,-26.5</points>
<connection>
<GID>1</GID>
<name>IN_4</name></connection>
<intersection>114.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>114.5,-37,142,-37</points>
<connection>
<GID>94</GID>
<name>IN_B_0</name></connection>
<intersection>114.5 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>114.5,6.5,119,6.5</points>
<connection>
<GID>487</GID>
<name>IN_4</name></connection>
<intersection>114.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>132,14.5,149.5,14.5</points>
<connection>
<GID>159</GID>
<name>IN_7</name></connection>
<intersection>149.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>149.5,12.5,149.5,25.5</points>
<intersection>12.5 17</intersection>
<intersection>14.5 2</intersection>
<intersection>25.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>149.5,25.5,151,25.5</points>
<connection>
<GID>428</GID>
<name>OUT_0</name></connection>
<intersection>149.5 9</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>149.5,12.5,167,12.5</points>
<connection>
<GID>423</GID>
<name>OUT_0</name></connection>
<intersection>149.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-27.5,113.5,5.5</points>
<intersection>-27.5 4</intersection>
<intersection>-9.5 1</intersection>
<intersection>-4.5 2</intersection>
<intersection>5.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-9.5,124.5,-9.5</points>
<connection>
<GID>196</GID>
<name>IN_3</name></connection>
<intersection>113.5 0</intersection>
<intersection>119 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-4.5,113.5,-4.5</points>
<connection>
<GID>194</GID>
<name>OUT_3</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>113.5,-27.5,124.5,-27.5</points>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>113.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>119,-18,119,-9.5</points>
<intersection>-18 6</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>119,-18,143,-18</points>
<connection>
<GID>87</GID>
<name>IN_B_3</name></connection>
<intersection>119 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>113.5,5.5,119,5.5</points>
<connection>
<GID>487</GID>
<name>IN_3</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-28.5,112.5,4.5</points>
<intersection>-28.5 4</intersection>
<intersection>-10.5 1</intersection>
<intersection>-3.5 2</intersection>
<intersection>4.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-10.5,124.5,-10.5</points>
<connection>
<GID>196</GID>
<name>IN_2</name></connection>
<intersection>112.5 0</intersection>
<intersection>119.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-3.5,112.5,-3.5</points>
<connection>
<GID>194</GID>
<name>OUT_2</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>112.5,-28.5,124.5,-28.5</points>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>112.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>119.5,-17,119.5,-10.5</points>
<intersection>-17 7</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>119.5,-17,143,-17</points>
<connection>
<GID>87</GID>
<name>IN_B_2</name></connection>
<intersection>119.5 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>112.5,4.5,119,4.5</points>
<connection>
<GID>487</GID>
<name>IN_2</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-5.5,139,0.5</points>
<intersection>-5.5 4</intersection>
<intersection>0 2</intersection>
<intersection>0.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>139,0,141,0</points>
<intersection>139 0</intersection>
<intersection>141 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>141,0,141,0.5</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>138,-5.5,139,-5.5</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>139,0.5,140,0.5</points>
<connection>
<GID>415</GID>
<name>clear</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-29.5,111.5,3.5</points>
<intersection>-29.5 4</intersection>
<intersection>-11.5 1</intersection>
<intersection>-2.5 2</intersection>
<intersection>3.5 10</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-11.5,124.5,-11.5</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>111.5 0</intersection>
<intersection>120 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-2.5,111.5,-2.5</points>
<connection>
<GID>194</GID>
<name>OUT_1</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111.5,-29.5,124.5,-29.5</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>111.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>120,-16,120,-11.5</points>
<intersection>-16 6</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>120,-16,143,-16</points>
<connection>
<GID>87</GID>
<name>IN_B_1</name></connection>
<intersection>120 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>111.5,3.5,119,3.5</points>
<connection>
<GID>487</GID>
<name>IN_1</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-5.5,144,-5.5</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<connection>
<GID>416</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-30.5,110.5,2.5</points>
<intersection>-30.5 4</intersection>
<intersection>-12.5 1</intersection>
<intersection>-1.5 2</intersection>
<intersection>2.5 13</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110.5,-12.5,124.5,-12.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>110.5 0</intersection>
<intersection>120.5 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-1.5,110.5,-1.5</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>110.5,-30.5,124.5,-30.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>120.5,-15,120.5,-12.5</points>
<intersection>-15 9</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>120.5,-15,143,-15</points>
<connection>
<GID>87</GID>
<name>IN_B_0</name></connection>
<intersection>120.5 8</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>110.5,2.5,119,2.5</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-5.5,134.5,13</points>
<intersection>-5.5 6</intersection>
<intersection>13 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>134.5,13,138,13</points>
<intersection>134.5 0</intersection>
<intersection>138 8</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>134.5,-5.5,136,-5.5</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>134.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>138,11.5,138,19.5</points>
<connection>
<GID>415</GID>
<name>load</name></connection>
<connection>
<GID>445</GID>
<name>OUT</name></connection>
<intersection>13 4</intersection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>152.5,-25.5,152.5,-25.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-6.5,140,-5.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,3.5,169,4</points>
<connection>
<GID>423</GID>
<name>ENABLE_0</name></connection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,3.5,169,3.5</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>169 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135.5,26.5,137,26.5</points>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<intersection>137 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>137,25.5,137,26.5</points>
<connection>
<GID>445</GID>
<name>IN_1</name></connection>
<intersection>26.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,26.5,131.5,26.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>161.5,-25.5,161.5,-20</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>-21 12</intersection>
<intersection>-20 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>161.5,-20,162.5,-20</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>161.5 2</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>161.5,-21,162.5,-21</points>
<connection>
<GID>88</GID>
<name>IN_2</name></connection>
<intersection>161.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,26.5,127.5,26.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>65,-19.5,67,-19.5</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<connection>
<GID>243</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,26.5,123.5,28.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-20.5,73,-20.5</points>
<connection>
<GID>247</GID>
<name>N_in0</name></connection>
<connection>
<GID>263</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>150,-40.5,171,-40.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<connection>
<GID>105</GID>
<name>IN_B_0</name></connection>
<intersection>151 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>151,-40.5,151,-34</points>
<intersection>-40.5 1</intersection>
<intersection>-34 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>151,-34,181,-34</points>
<connection>
<GID>95</GID>
<name>IN_B_0</name></connection>
<intersection>151 6</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>150,-42.5,171,-42.5</points>
<connection>
<GID>94</GID>
<name>OUT_2</name></connection>
<connection>
<GID>105</GID>
<name>IN_B_2</name></connection>
<intersection>152 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>152,-42.5,152,-36</points>
<intersection>-42.5 1</intersection>
<intersection>-36 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>152,-36,181,-36</points>
<connection>
<GID>95</GID>
<name>IN_B_2</name></connection>
<intersection>152 6</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>150,-41.5,171,-41.5</points>
<connection>
<GID>94</GID>
<name>OUT_1</name></connection>
<connection>
<GID>105</GID>
<name>IN_B_1</name></connection>
<intersection>151.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>151.5,-41.5,151.5,-35</points>
<intersection>-41.5 1</intersection>
<intersection>-35 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>151.5,-35,181,-35</points>
<connection>
<GID>95</GID>
<name>IN_B_1</name></connection>
<intersection>151.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>150,-43.5,171,-43.5</points>
<connection>
<GID>94</GID>
<name>OUT_3</name></connection>
<connection>
<GID>105</GID>
<name>IN_B_3</name></connection>
<intersection>152.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>152.5,-43.5,152.5,-37</points>
<intersection>-43.5 1</intersection>
<intersection>-37 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>152.5,-37,181,-37</points>
<connection>
<GID>95</GID>
<name>IN_B_3</name></connection>
<intersection>152.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-26,66.5,-21.5</points>
<intersection>-26 5</intersection>
<intersection>-21.5 15</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>62.5,-26,76,-26</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>66.5,-21.5,67,-21.5</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,94,237.5,94</points>
<connection>
<GID>446</GID>
<name>OUT</name></connection>
<connection>
<GID>470</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,96,231.5,96</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<connection>
<GID>447</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51,-24.5,52.5,-24.5</points>
<connection>
<GID>237</GID>
<name>clear</name></connection>
<connection>
<GID>237</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,89,231.5,92</points>
<connection>
<GID>524</GID>
<name>OUT</name></connection>
<connection>
<GID>446</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>17</ID>
<points>121,15,121,36.5</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>22.5 19</intersection>
<intersection>32.5 23</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>121,22.5,133.5,22.5</points>
<intersection>121 17</intersection>
<intersection>133.5 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>133.5,12.5,133.5,22.5</points>
<connection>
<GID>159</GID>
<name>ENABLE_0</name></connection>
<intersection>22.5 19</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>121,32.5,123.5,32.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>121 17</intersection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,93,231.5,94</points>
<connection>
<GID>448</GID>
<name>OUT</name></connection>
<connection>
<GID>446</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>180,-47.5,180,-42</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>-43 7</intersection>
<intersection>-42 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>180,-43,181,-43</points>
<connection>
<GID>95</GID>
<name>IN_2</name></connection>
<intersection>180 2</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>180,-42,181,-42</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>180 2</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-34,145,-28</points>
<connection>
<GID>94</GID>
<name>carry_in</name></connection>
<intersection>-34 1</intersection>
<intersection>-28 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-34,162.5,-34</points>
<intersection>145 0</intersection>
<intersection>162.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>162.5,-34,162.5,-31.5</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-28,146,-28</points>
<connection>
<GID>87</GID>
<name>carry_out</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,31,227,33.5</points>
<intersection>31 2</intersection>
<intersection>33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226,33.5,227,33.5</points>
<connection>
<GID>442</GID>
<name>OUT</name></connection>
<intersection>227 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,31,228.5,31</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>227 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-21,177,12.5</points>
<intersection>-21 2</intersection>
<intersection>-18.5 1</intersection>
<intersection>12.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170.5,-18.5,177,-18.5</points>
<connection>
<GID>88</GID>
<name>OUT_3</name></connection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,-21,217,-21</points>
<connection>
<GID>108</GID>
<name>IN_3</name></connection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>171,12.5,177,12.5</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<intersection>177 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-22,217,-22</points>
<connection>
<GID>108</GID>
<name>IN_2</name></connection>
<intersection>170 9</intersection>
<intersection>175.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>175.5,-22,175.5,11.5</points>
<intersection>-22 1</intersection>
<intersection>11.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>171,11.5,175.5,11.5</points>
<connection>
<GID>423</GID>
<name>IN_1</name></connection>
<intersection>175.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>170,-22,170,-17.5</points>
<intersection>-22 1</intersection>
<intersection>-17.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>170,-17.5,170.5,-17.5</points>
<connection>
<GID>88</GID>
<name>OUT_2</name></connection>
<intersection>170 9</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-23,217,-23</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>177 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>177,-23,177,-16.5</points>
<intersection>-23 1</intersection>
<intersection>-16.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>170.5,-16.5,177,-16.5</points>
<connection>
<GID>88</GID>
<name>OUT_1</name></connection>
<intersection>174 5</intersection>
<intersection>177 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>174,-16.5,174,10.5</points>
<intersection>-16.5 4</intersection>
<intersection>10.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>171,10.5,174,10.5</points>
<connection>
<GID>423</GID>
<name>IN_2</name></connection>
<intersection>174 5</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-14.5,53.5,-12</points>
<connection>
<GID>237</GID>
<name>load</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-12,85.5,-12</points>
<intersection>53.5 0</intersection>
<intersection>84 16</intersection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-12,85.5,8</points>
<intersection>-12 1</intersection>
<intersection>-9.5 5</intersection>
<intersection>8 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>78.5,8,85.5,8</points>
<intersection>78.5 7</intersection>
<intersection>85.5 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>78.5,-9.5,85.5,-9.5</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>78.5 8</intersection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>78.5,3.5,78.5,8</points>
<connection>
<GID>107</GID>
<name>load</name></connection>
<intersection>8 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>78.5,-9.5,78.5,-7.5</points>
<connection>
<GID>107</GID>
<name>clock</name></connection>
<intersection>-9.5 5</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>84,-15,84,-12</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-24,177,-15.5</points>
<intersection>-24 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170.5,-15.5,177,-15.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<intersection>172 3</intersection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,-24,217,-24</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>172,-15.5,172,9.5</points>
<intersection>-15.5 1</intersection>
<intersection>9.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>171,9.5,172,9.5</points>
<connection>
<GID>423</GID>
<name>IN_3</name></connection>
<intersection>172 3</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-11,101.5,-9</points>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<connection>
<GID>197</GID>
<name>shift_left</name></connection></vsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>158.5,-32,160.5,-32</points>
<intersection>158.5 6</intersection>
<intersection>160.5 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>158.5,-32,158.5,-31.5</points>
<connection>
<GID>89</GID>
<name>A_less_B</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>160.5,-32,160.5,-31.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-26,80,-26</points>
<connection>
<GID>291</GID>
<name>OUT_0</name></connection>
<connection>
<GID>292</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-26,103.5,28</points>
<intersection>-26 8</intersection>
<intersection>-21 5</intersection>
<intersection>-8 6</intersection>
<intersection>28 13</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>100.5,-21,103.5,-21</points>
<connection>
<GID>197</GID>
<name>clock</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>100.5,-8,103.5,-8</points>
<connection>
<GID>194</GID>
<name>clock</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>92,-26,103.5,-26</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>103.5,28,105,28</points>
<connection>
<GID>155</GID>
<name>clock</name></connection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-26,88,-26</points>
<connection>
<GID>293</GID>
<name>OUT_0</name></connection>
<connection>
<GID>294</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-26,84,-26</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<connection>
<GID>293</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189,-37.5,197,-37.5</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>190 10</intersection>
<intersection>197 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>197,-37.5,197,-31</points>
<intersection>-37.5 1</intersection>
<intersection>-31 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>197,-31,210,-31</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>197 3</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>190,-37.5,190,5.5</points>
<intersection>-37.5 1</intersection>
<intersection>5.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>171,5.5,190,5.5</points>
<connection>
<GID>423</GID>
<name>IN_7</name></connection>
<intersection>190 10</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189,-38.5,197,-38.5</points>
<connection>
<GID>95</GID>
<name>OUT_1</name></connection>
<intersection>191.5 8</intersection>
<intersection>197 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>197,-38.5,197,-30</points>
<intersection>-38.5 1</intersection>
<intersection>-30 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>197,-30,210,-30</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>197 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>191.5,-38.5,191.5,6.5</points>
<intersection>-38.5 1</intersection>
<intersection>6.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>171,6.5,191.5,6.5</points>
<connection>
<GID>423</GID>
<name>IN_6</name></connection>
<intersection>191.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189,-39.5,197,-39.5</points>
<connection>
<GID>95</GID>
<name>OUT_2</name></connection>
<intersection>192.5 9</intersection>
<intersection>197 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>197,-39.5,197,-29</points>
<intersection>-39.5 1</intersection>
<intersection>-29 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>197,-29,210,-29</points>
<connection>
<GID>110</GID>
<name>IN_2</name></connection>
<intersection>197 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>192.5,-39.5,192.5,7.5</points>
<intersection>-39.5 1</intersection>
<intersection>7.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>171,7.5,192.5,7.5</points>
<connection>
<GID>423</GID>
<name>IN_5</name></connection>
<intersection>192.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189,-40.5,197,-40.5</points>
<connection>
<GID>95</GID>
<name>OUT_3</name></connection>
<intersection>193.5 8</intersection>
<intersection>197 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>197,-40.5,197,-28</points>
<intersection>-40.5 1</intersection>
<intersection>-28 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>197,-28,210,-28</points>
<connection>
<GID>110</GID>
<name>IN_3</name></connection>
<intersection>197 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>193.5,-40.5,193.5,8.5</points>
<intersection>-40.5 1</intersection>
<intersection>8.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>171,8.5,193.5,8.5</points>
<connection>
<GID>423</GID>
<name>IN_4</name></connection>
<intersection>193.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>226,29,228.5,29</points>
<connection>
<GID>460</GID>
<name>OUT</name></connection>
<connection>
<GID>459</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>630</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226,24.5,226,27</points>
<intersection>24.5 2</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226,27,228.5,27</points>
<connection>
<GID>459</GID>
<name>IN_2</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,24.5,226,24.5</points>
<connection>
<GID>461</GID>
<name>OUT</name></connection>
<intersection>226 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165.5,-46.5,165.5,-25</points>
<connection>
<GID>88</GID>
<name>carry_out</name></connection>
<intersection>-46.5 25</intersection>
<intersection>-26 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>165.5,-26,184,-26</points>
<intersection>165.5 0</intersection>
<intersection>184 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>184,-31,184,-26</points>
<connection>
<GID>95</GID>
<name>carry_in</name></connection>
<intersection>-26 3</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>165,-46.5,165.5,-46.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>631</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,19,227,25</points>
<intersection>19 2</intersection>
<intersection>25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227,25,228.5,25</points>
<connection>
<GID>459</GID>
<name>IN_3</name></connection>
<intersection>227 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>226,19,227,19</points>
<connection>
<GID>450</GID>
<name>OUT</name></connection>
<intersection>227 0</intersection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,19,220,19</points>
<connection>
<GID>450</GID>
<name>IN_1</name></connection>
<connection>
<GID>467</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>171,-47.5,171,-47.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<connection>
<GID>112</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>241.5,126.5,241.5,126.5</points>
<connection>
<GID>486</GID>
<name>OUT</name></connection>
<connection>
<GID>489</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-30.5,141.5,-22</points>
<intersection>-30.5 2</intersection>
<intersection>-22 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-30.5,141.5,-30.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>141.5,-22,143,-22</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,119.5,234.5,123.5</points>
<connection>
<GID>486</GID>
<name>IN_3</name></connection>
<intersection>119.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>234,119.5,234.5,119.5</points>
<connection>
<GID>484</GID>
<name>OUT</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-29.5,142,-23</points>
<intersection>-29.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-23,143,-23</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-29.5,142,-29.5</points>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,123.5,234,125.5</points>
<connection>
<GID>483</GID>
<name>OUT</name></connection>
<intersection>125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,125.5,234.5,125.5</points>
<connection>
<GID>486</GID>
<name>IN_2</name></connection>
<intersection>234 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-28.5,142.5,-24</points>
<intersection>-28.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142.5,-24,143,-24</points>
<connection>
<GID>87</GID>
<name>IN_2</name></connection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-28.5,142.5,-28.5</points>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<intersection>142.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,79,177,130.5</points>
<intersection>79 2</intersection>
<intersection>110.5 6</intersection>
<intersection>130.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,130.5,234.5,130.5</points>
<intersection>177 0</intersection>
<intersection>234.5 23</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>175.5,79,230,79</points>
<intersection>175.5 35</intersection>
<intersection>177 0</intersection>
<intersection>230 21</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>177,110.5,245.5,110.5</points>
<intersection>177 0</intersection>
<intersection>245.5 24</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>230,76,230,79</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>79 2</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>234.5,129.5,234.5,130.5</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>130.5 1</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>245.5,110,245.5,110.5</points>
<connection>
<GID>464</GID>
<name>IN_1</name></connection>
<intersection>110.5 6</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>175.5,68.5,175.5,79</points>
<intersection>68.5 36</intersection>
<intersection>79 2</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>172,68.5,175.5,68.5</points>
<connection>
<GID>656</GID>
<name>N_in1</name></connection>
<intersection>175.5 35</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-27.5,143,-25</points>
<connection>
<GID>87</GID>
<name>IN_3</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-27.5,143,-27.5</points>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,122.5,228,122.5</points>
<connection>
<GID>483</GID>
<name>IN_1</name></connection>
<connection>
<GID>490</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-44,138,-26.5</points>
<intersection>-44 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-26.5,138,-26.5</points>
<connection>
<GID>1</GID>
<name>OUT_4</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-44,142,-44</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,118.5,228,118.5</points>
<connection>
<GID>520</GID>
<name>OUT_0</name></connection>
<connection>
<GID>484</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-45,138.5,-25.5</points>
<intersection>-45 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-25.5,138.5,-25.5</points>
<connection>
<GID>1</GID>
<name>OUT_5</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,-45,142,-45</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,71,219,71</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>177 52</intersection>
<intersection>189 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>189,17,189,126.5</points>
<intersection>17 47</intersection>
<intersection>23.5 42</intersection>
<intersection>32.5 22</intersection>
<intersection>40.5 51</intersection>
<intersection>51.5 30</intersection>
<intersection>55.5 18</intersection>
<intersection>71 1</intersection>
<intersection>88 37</intersection>
<intersection>103 28</intersection>
<intersection>107 38</intersection>
<intersection>118.5 8</intersection>
<intersection>126.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>189,126.5,228,126.5</points>
<connection>
<GID>523</GID>
<name>IN_1</name></connection>
<intersection>189 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>189,118.5,218,118.5</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<intersection>189 5</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>189,55.5,224.5,55.5</points>
<connection>
<GID>455</GID>
<name>IN_1</name></connection>
<intersection>189 5</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>189,32.5,220,32.5</points>
<connection>
<GID>442</GID>
<name>IN_1</name></connection>
<intersection>189 5</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>189,103,239.5,103</points>
<connection>
<GID>466</GID>
<name>IN_1</name></connection>
<intersection>189 5</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>189,51.5,220.5,51.5</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>189 5</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>189,88,225.5,88</points>
<connection>
<GID>524</GID>
<name>IN_1</name></connection>
<intersection>189 5</intersection>
<intersection>193 44</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>189,107,239.5,107</points>
<connection>
<GID>465</GID>
<name>IN_1</name></connection>
<intersection>189 5</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>189,23.5,213.5,23.5</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>189 5</intersection></hsegment>
<vsegment>
<ID>44</ID>
<points>193,88,193,92</points>
<intersection>88 37</intersection>
<intersection>92 45</intersection></vsegment>
<hsegment>
<ID>45</ID>
<points>193,92,225.5,92</points>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<intersection>193 44</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>189,17,220,17</points>
<connection>
<GID>450</GID>
<name>IN_2</name></connection>
<intersection>189 5</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>189,40.5,228,40.5</points>
<connection>
<GID>457</GID>
<name>IN_2</name></connection>
<intersection>189 5</intersection></hsegment>
<vsegment>
<ID>52</ID>
<points>177,64.5,177,71</points>
<intersection>64.5 53</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>172,64.5,177,64.5</points>
<connection>
<GID>638</GID>
<name>N_in1</name></connection>
<intersection>177 52</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-46,139,-24.5</points>
<intersection>-46 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-24.5,139,-24.5</points>
<connection>
<GID>1</GID>
<name>OUT_6</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139,-46,142,-46</points>
<connection>
<GID>94</GID>
<name>IN_2</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180,21,180,124.5</points>
<intersection>21 41</intersection>
<intersection>30 37</intersection>
<intersection>34.5 17</intersection>
<intersection>42.5 45</intersection>
<intersection>57.5 30</intersection>
<intersection>67 47</intersection>
<intersection>69 15</intersection>
<intersection>77 5</intersection>
<intersection>96 39</intersection>
<intersection>105 25</intersection>
<intersection>109 11</intersection>
<intersection>120.5 1</intersection>
<intersection>124.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180,120.5,228,120.5</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>180,124.5,228,124.5</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>180,77,219,77</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>180,109,239.5,109</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>180,69,223,69</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>180,34.5,220,34.5</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>180,105,239.5,105</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>180,57.5,224.5,57.5</points>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>180,30,208,30</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>180,96,227.5,96</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>180,21,220,21</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>180,42.5,228,42.5</points>
<connection>
<GID>457</GID>
<name>IN_1</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>172,67,180,67</points>
<connection>
<GID>655</GID>
<name>N_in1</name></connection>
<intersection>180 0</intersection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-47,139.5,-23.5</points>
<intersection>-47 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-23.5,139.5,-23.5</points>
<connection>
<GID>1</GID>
<name>OUT_7</name></connection>
<intersection>139.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139.5,-47,142,-47</points>
<connection>
<GID>94</GID>
<name>IN_3</name></connection>
<intersection>139.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,19,185,128.5</points>
<intersection>19 33</intersection>
<intersection>25.5 28</intersection>
<intersection>28 18</intersection>
<intersection>44.5 16</intersection>
<intersection>53.5 25</intersection>
<intersection>67 12</intersection>
<intersection>73 1</intersection>
<intersection>75 8</intersection>
<intersection>90 26</intersection>
<intersection>94 31</intersection>
<intersection>112 22</intersection>
<intersection>122.5 2</intersection>
<intersection>128.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178,73,223,73</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>178 36</intersection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,122.5,224,122.5</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>185,128.5,228,128.5</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>185,75,223,75</points>
<connection>
<GID>526</GID>
<name>IN_1</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>185,67,219,67</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>185,44.5,224,44.5</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>185,28,220,28</points>
<connection>
<GID>460</GID>
<name>IN_1</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>185,112,245.5,112</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>185,53.5,224.5,53.5</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>185,90,225.5,90</points>
<connection>
<GID>524</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>185,25.5,219.5,25.5</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>185,94,225.5,94</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>185,19,216,19</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>178,65.5,178,73</points>
<intersection>65.5 37</intersection>
<intersection>73 1</intersection></vsegment>
<hsegment>
<ID>37</ID>
<points>172,65.5,178,65.5</points>
<connection>
<GID>654</GID>
<name>N_in1</name></connection>
<intersection>178 36</intersection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234,127.5,234.5,127.5</points>
<connection>
<GID>523</GID>
<name>OUT</name></connection>
<connection>
<GID>486</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,74,229,76</points>
<connection>
<GID>526</GID>
<name>OUT</name></connection>
<intersection>74 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>229,74,230,74</points>
<connection>
<GID>525</GID>
<name>IN_1</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-25,93,-8</points>
<intersection>-25 4</intersection>
<intersection>-8 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>93,-8,99.5,-8</points>
<connection>
<GID>194</GID>
<name>clear</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>93,-25,99.5,-25</points>
<intersection>93 0</intersection>
<intersection>99.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>99.5,-28,99.5,-21</points>
<connection>
<GID>197</GID>
<name>clear</name></connection>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>-25 4</intersection></vsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>229,72,230,72</points>
<connection>
<GID>527</GID>
<name>OUT</name></connection>
<connection>
<GID>525</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>100.5,-34,100.5,-34</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,68,229.5,70</points>
<intersection>68 1</intersection>
<intersection>70 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229,68,229.5,68</points>
<connection>
<GID>468</GID>
<name>OUT</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>229.5,70,230,70</points>
<connection>
<GID>525</GID>
<name>IN_3</name></connection>
<intersection>229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>98.5,-34,98.5,-34</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<connection>
<GID>116</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223,77,223,77</points>
<connection>
<GID>449</GID>
<name>OUT_0</name></connection>
<connection>
<GID>526</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-33,127.5,-32.5</points>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<connection>
<GID>118</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223,71,223,71</points>
<connection>
<GID>451</GID>
<name>OUT_0</name></connection>
<connection>
<GID>527</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-41,132,-32.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-41 5</intersection>
<intersection>-32.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>129.5,-32.5,132,-32.5</points>
<connection>
<GID>1</GID>
<name>clear</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>128.5,-41,132,-41</points>
<intersection>128.5 6</intersection>
<intersection>132 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>128.5,-41,128.5,-39</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>-41 5</intersection></vsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223,67,223,67</points>
<connection>
<GID>452</GID>
<name>OUT_0</name></connection>
<connection>
<GID>468</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,73,237,73</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<connection>
<GID>525</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,55,236.5,55</points>
<connection>
<GID>453</GID>
<name>OUT</name></connection>
<connection>
<GID>474</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,52.5,230.5,54</points>
<connection>
<GID>454</GID>
<name>OUT</name></connection>
<connection>
<GID>453</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,56,230.5,56.5</points>
<connection>
<GID>455</GID>
<name>OUT</name></connection>
<connection>
<GID>453</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224.5,51.5,224.5,51.5</points>
<connection>
<GID>454</GID>
<name>IN_1</name></connection>
<connection>
<GID>456</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,42.5,234,42.5</points>
<connection>
<GID>457</GID>
<name>OUT</name></connection>
<connection>
<GID>482</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,44.5,228,44.5</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<connection>
<GID>458</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235.5,28,236.5,28</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<connection>
<GID>459</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212,30,220,30</points>
<connection>
<GID>462</GID>
<name>OUT_0</name></connection>
<connection>
<GID>460</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>658</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217.5,23.5,219.5,23.5</points>
<connection>
<GID>463</GID>
<name>OUT_0</name></connection>
<connection>
<GID>461</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>659</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>252.5,109,252.5,109</points>
<connection>
<GID>464</GID>
<name>OUT</name></connection>
<connection>
<GID>469</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>660</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,108,245.5,108</points>
<connection>
<GID>464</GID>
<name>IN_2</name></connection>
<connection>
<GID>465</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,104,245.5,106</points>
<connection>
<GID>466</GID>
<name>OUT</name></connection>
<connection>
<GID>464</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336,96,336,96</points>
<connection>
<GID>529</GID>
<name>OUT</name></connection>
<connection>
<GID>553</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,98,330,98</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<connection>
<GID>530</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>664</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,91,330,94</points>
<connection>
<GID>566</GID>
<name>OUT</name></connection>
<connection>
<GID>529</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>665</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,95,330,96</points>
<connection>
<GID>531</GID>
<name>OUT</name></connection>
<connection>
<GID>529</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325.5,33,325.5,37.5</points>
<intersection>33 2</intersection>
<intersection>37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>324,37.5,325.5,37.5</points>
<connection>
<GID>528</GID>
<name>OUT</name></connection>
<intersection>325.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>325.5,33,327,33</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<intersection>325.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>667</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>324.5,31,327,31</points>
<connection>
<GID>543</GID>
<name>OUT</name></connection>
<connection>
<GID>542</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>668</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>324.5,26.5,324.5,29</points>
<intersection>26.5 2</intersection>
<intersection>29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>324.5,29,327,29</points>
<connection>
<GID>542</GID>
<name>IN_2</name></connection>
<intersection>324.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>324,26.5,324.5,26.5</points>
<connection>
<GID>544</GID>
<name>OUT</name></connection>
<intersection>324.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325.5,21,325.5,27</points>
<intersection>21 2</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>325.5,27,327,27</points>
<connection>
<GID>542</GID>
<name>IN_3</name></connection>
<intersection>325.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>324.5,21,325.5,21</points>
<connection>
<GID>533</GID>
<name>OUT</name></connection>
<intersection>325.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318.5,21,318.5,21</points>
<connection>
<GID>533</GID>
<name>IN_1</name></connection>
<connection>
<GID>550</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,9.5,125,10.5</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,9.5,135,9.5</points>
<connection>
<GID>415</GID>
<name>IN_7</name></connection>
<connection>
<GID>487</GID>
<name>OUT_7</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>340,128.5,340,128.5</points>
<connection>
<GID>561</GID>
<name>OUT</name></connection>
<connection>
<GID>562</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,121.5,333,125.5</points>
<connection>
<GID>561</GID>
<name>IN_3</name></connection>
<intersection>121.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>332.5,121.5,333,121.5</points>
<connection>
<GID>559</GID>
<name>OUT</name></connection>
<intersection>333 0</intersection></hsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332.5,125.5,332.5,127.5</points>
<connection>
<GID>558</GID>
<name>OUT</name></connection>
<intersection>127.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>332.5,127.5,333,127.5</points>
<connection>
<GID>561</GID>
<name>IN_2</name></connection>
<intersection>332.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,8.5,135,8.5</points>
<connection>
<GID>415</GID>
<name>IN_6</name></connection>
<connection>
<GID>487</GID>
<name>OUT_6</name></connection>
<intersection>126 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>126,8.5,126,10.5</points>
<connection>
<GID>159</GID>
<name>OUT_1</name></connection>
<intersection>8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275.5,81,275.5,132.5</points>
<intersection>81 2</intersection>
<intersection>112.5 6</intersection>
<intersection>132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275.5,132.5,333,132.5</points>
<intersection>275.5 0</intersection>
<intersection>333 23</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>273,81,328.5,81</points>
<intersection>273 29</intersection>
<intersection>275.5 0</intersection>
<intersection>328.5 21</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>275.5,112.5,344,112.5</points>
<intersection>275.5 0</intersection>
<intersection>344 24</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>328.5,78,328.5,81</points>
<connection>
<GID>567</GID>
<name>IN_0</name></connection>
<intersection>81 2</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>333,131.5,333,132.5</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>132.5 1</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>344,112,344,112.5</points>
<connection>
<GID>547</GID>
<name>IN_1</name></connection>
<intersection>112.5 6</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>273,67.5,273,81</points>
<intersection>67.5 34</intersection>
<intersection>81 2</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>269.5,67.5,273,67.5</points>
<connection>
<GID>664</GID>
<name>N_in1</name></connection>
<intersection>273 29</intersection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,7.5,135,7.5</points>
<connection>
<GID>415</GID>
<name>IN_5</name></connection>
<connection>
<GID>487</GID>
<name>OUT_5</name></connection>
<intersection>127 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>127,7.5,127,10.5</points>
<connection>
<GID>159</GID>
<name>OUT_2</name></connection>
<intersection>7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326.5,124.5,326.5,124.5</points>
<connection>
<GID>558</GID>
<name>IN_1</name></connection>
<connection>
<GID>563</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>320.5,120.5,326.5,120.5</points>
<connection>
<GID>564</GID>
<name>OUT_0</name></connection>
<connection>
<GID>559</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>677</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>275,73,317.5,73</points>
<connection>
<GID>534</GID>
<name>IN_0</name></connection>
<intersection>275 50</intersection>
<intersection>287.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>287.5,19,287.5,128.5</points>
<intersection>19 47</intersection>
<intersection>25.5 42</intersection>
<intersection>36.5 40</intersection>
<intersection>42.5 22</intersection>
<intersection>53.5 30</intersection>
<intersection>57.5 18</intersection>
<intersection>73 1</intersection>
<intersection>90 37</intersection>
<intersection>105 28</intersection>
<intersection>109 38</intersection>
<intersection>120.5 8</intersection>
<intersection>128.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>287.5,128.5,326.5,128.5</points>
<connection>
<GID>565</GID>
<name>IN_1</name></connection>
<intersection>287.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>287.5,120.5,316.5,120.5</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>287.5 5</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>287.5,57.5,323,57.5</points>
<connection>
<GID>538</GID>
<name>IN_1</name></connection>
<intersection>287.5 5</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>287.5,42.5,326.5,42.5</points>
<connection>
<GID>540</GID>
<name>IN_2</name></connection>
<intersection>287.5 5</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>287.5,105,338,105</points>
<connection>
<GID>549</GID>
<name>IN_1</name></connection>
<intersection>287.5 5</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>287.5,53.5,319,53.5</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>287.5 5</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>287.5,90,324,90</points>
<connection>
<GID>566</GID>
<name>IN_1</name></connection>
<intersection>287.5 5</intersection>
<intersection>291.5 44</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>287.5,109,338,109</points>
<connection>
<GID>548</GID>
<name>IN_1</name></connection>
<intersection>287.5 5</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>287.5,36.5,318,36.5</points>
<connection>
<GID>528</GID>
<name>IN_1</name></connection>
<intersection>287.5 5</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>287.5,25.5,312,25.5</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>287.5 5</intersection></hsegment>
<vsegment>
<ID>44</ID>
<points>291.5,90,291.5,94</points>
<intersection>90 37</intersection>
<intersection>94 45</intersection></vsegment>
<hsegment>
<ID>45</ID>
<points>291.5,94,324,94</points>
<connection>
<GID>531</GID>
<name>IN_1</name></connection>
<intersection>291.5 44</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>287.5,19,318.5,19</points>
<connection>
<GID>533</GID>
<name>IN_2</name></connection>
<intersection>287.5 5</intersection></hsegment>
<vsegment>
<ID>50</ID>
<points>275,63.5,275,73</points>
<intersection>63.5 51</intersection>
<intersection>73 1</intersection></vsegment>
<hsegment>
<ID>51</ID>
<points>269.5,63.5,275,63.5</points>
<connection>
<GID>661</GID>
<name>N_in1</name></connection>
<intersection>275 50</intersection></hsegment></shape></wire>
<wire>
<ID>678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278.5,23,278.5,126.5</points>
<intersection>23 41</intersection>
<intersection>32 37</intersection>
<intersection>38.5 35</intersection>
<intersection>44.5 17</intersection>
<intersection>59.5 30</intersection>
<intersection>66 45</intersection>
<intersection>71 15</intersection>
<intersection>79 5</intersection>
<intersection>98 39</intersection>
<intersection>107 25</intersection>
<intersection>111 11</intersection>
<intersection>122.5 1</intersection>
<intersection>126.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278.5,122.5,326.5,122.5</points>
<connection>
<GID>559</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>278.5,126.5,326.5,126.5</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>278.5,79,317.5,79</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>278.5,111,338,111</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>278.5,71,321.5,71</points>
<connection>
<GID>551</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>278.5,44.5,326.5,44.5</points>
<connection>
<GID>540</GID>
<name>IN_1</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>278.5,107,338,107</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>278.5,59.5,323,59.5</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>278.5,38.5,318,38.5</points>
<connection>
<GID>528</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>278.5,32,306.5,32</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>278.5,98,326,98</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>278.5,23,318.5,23</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>269.5,66,278.5,66</points>
<connection>
<GID>663</GID>
<name>N_in1</name></connection>
<intersection>278.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>283.5,21,283.5,130.5</points>
<intersection>21 33</intersection>
<intersection>27.5 28</intersection>
<intersection>30 18</intersection>
<intersection>46.5 16</intersection>
<intersection>55.5 25</intersection>
<intersection>69 12</intersection>
<intersection>75 1</intersection>
<intersection>77 8</intersection>
<intersection>92 26</intersection>
<intersection>96 31</intersection>
<intersection>114 22</intersection>
<intersection>124.5 2</intersection>
<intersection>130.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,75,321.5,75</points>
<connection>
<GID>569</GID>
<name>IN_0</name></connection>
<intersection>274 36</intersection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>283.5,124.5,322.5,124.5</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>283.5,130.5,326.5,130.5</points>
<connection>
<GID>565</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>283.5,77,321.5,77</points>
<connection>
<GID>568</GID>
<name>IN_1</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>283.5,69,317.5,69</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>283.5,46.5,322.5,46.5</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>283.5,30,318.5,30</points>
<connection>
<GID>543</GID>
<name>IN_1</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>283.5,114,344,114</points>
<connection>
<GID>547</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>283.5,55.5,323,55.5</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>283.5,92,324,92</points>
<connection>
<GID>566</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>283.5,27.5,318,27.5</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>283.5,96,324,96</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>283.5,21,314.5,21</points>
<connection>
<GID>550</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>274,64.5,274,75</points>
<intersection>64.5 37</intersection>
<intersection>75 1</intersection></vsegment>
<hsegment>
<ID>37</ID>
<points>269.5,64.5,274,64.5</points>
<connection>
<GID>662</GID>
<name>N_in1</name></connection>
<intersection>274 36</intersection></hsegment></shape></wire>
<wire>
<ID>680</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>332.5,129.5,333,129.5</points>
<connection>
<GID>565</GID>
<name>OUT</name></connection>
<connection>
<GID>561</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327.5,76,327.5,78</points>
<connection>
<GID>568</GID>
<name>OUT</name></connection>
<intersection>76 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>327.5,76,328.5,76</points>
<connection>
<GID>567</GID>
<name>IN_1</name></connection>
<intersection>327.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>682</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>327.5,74,328.5,74</points>
<connection>
<GID>569</GID>
<name>OUT</name></connection>
<connection>
<GID>567</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328,70,328,72</points>
<intersection>70 1</intersection>
<intersection>72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>327.5,70,328,70</points>
<connection>
<GID>551</GID>
<name>OUT</name></connection>
<intersection>328 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>328,72,328.5,72</points>
<connection>
<GID>567</GID>
<name>IN_3</name></connection>
<intersection>328 0</intersection></hsegment></shape></wire>
<wire>
<ID>684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321.5,79,321.5,79</points>
<connection>
<GID>532</GID>
<name>OUT_0</name></connection>
<connection>
<GID>568</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321.5,73,321.5,73</points>
<connection>
<GID>534</GID>
<name>OUT_0</name></connection>
<connection>
<GID>569</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>686</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321.5,69,321.5,69</points>
<connection>
<GID>535</GID>
<name>OUT_0</name></connection>
<connection>
<GID>551</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>687</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335.5,75,335.5,75</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<connection>
<GID>567</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335,57,335,57</points>
<connection>
<GID>536</GID>
<name>OUT</name></connection>
<connection>
<GID>555</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329,54.5,329,56</points>
<connection>
<GID>537</GID>
<name>OUT</name></connection>
<connection>
<GID>536</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329,58,329,58.5</points>
<connection>
<GID>538</GID>
<name>OUT</name></connection>
<connection>
<GID>536</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323,53.5,323,53.5</points>
<connection>
<GID>537</GID>
<name>IN_1</name></connection>
<connection>
<GID>539</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332.5,44.5,332.5,44.5</points>
<connection>
<GID>540</GID>
<name>OUT</name></connection>
<connection>
<GID>557</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326.5,46.5,326.5,46.5</points>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<connection>
<GID>541</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>334,30,335,30</points>
<connection>
<GID>542</GID>
<name>OUT</name></connection>
<connection>
<GID>556</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>310.5,32,318.5,32</points>
<connection>
<GID>545</GID>
<name>OUT_0</name></connection>
<connection>
<GID>543</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>316,25.5,318,25.5</points>
<connection>
<GID>546</GID>
<name>OUT_0</name></connection>
<connection>
<GID>544</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351,111,351,111</points>
<connection>
<GID>547</GID>
<name>OUT</name></connection>
<connection>
<GID>552</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344,110,344,110</points>
<connection>
<GID>547</GID>
<name>IN_2</name></connection>
<connection>
<GID>548</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344,106,344,108</points>
<connection>
<GID>549</GID>
<name>OUT</name></connection>
<connection>
<GID>547</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>722</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,43,85,43</points>
<connection>
<GID>614</GID>
<name>OUT_0</name></connection>
<connection>
<GID>621</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>723</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,43,89,43</points>
<connection>
<GID>613</GID>
<name>OUT_0</name></connection>
<connection>
<GID>622</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>724</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,43,93,43</points>
<connection>
<GID>612</GID>
<name>OUT_0</name></connection>
<connection>
<GID>623</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>725</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,35.5,85,35.5</points>
<connection>
<GID>617</GID>
<name>OUT_0</name></connection>
<connection>
<GID>624</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>726</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,35.5,89,35.5</points>
<connection>
<GID>616</GID>
<name>OUT_0</name></connection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89,35.5,89,35.5</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>727</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>93,35.5,93,35.5</points>
<connection>
<GID>615</GID>
<name>OUT_0</name></connection>
<connection>
<GID>626</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>728</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,28,85,28</points>
<connection>
<GID>620</GID>
<name>OUT_0</name></connection>
<connection>
<GID>627</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>729</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,28,89,28</points>
<connection>
<GID>619</GID>
<name>OUT_0</name></connection>
<connection>
<GID>628</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,28,93,28</points>
<connection>
<GID>618</GID>
<name>OUT_0</name></connection>
<connection>
<GID>629</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,20.5,89,20.5</points>
<connection>
<GID>611</GID>
<name>OUT_0</name></connection>
<connection>
<GID>630</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,42.5,99,42.5</points>
<connection>
<GID>631</GID>
<name>OUT_0</name></connection>
<connection>
<GID>632</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>96,42.5,96,43</points>
<connection>
<GID>633</GID>
<name>OUT_0</name></connection>
<connection>
<GID>634</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,42.5,102,42.5</points>
<connection>
<GID>635</GID>
<name>OUT_0</name></connection>
<connection>
<GID>636</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>759</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,11,121,11</points>
<connection>
<GID>487</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>519</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>760</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143.5,9.5,143.5,68.5</points>
<intersection>9.5 1</intersection>
<intersection>68.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,9.5,143.5,9.5</points>
<connection>
<GID>415</GID>
<name>OUT_7</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,68.5,170,68.5</points>
<connection>
<GID>656</GID>
<name>N_in0</name></connection>
<intersection>143.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>761</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,8.5,144,67</points>
<intersection>8.5 1</intersection>
<intersection>67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,8.5,144,8.5</points>
<connection>
<GID>415</GID>
<name>OUT_6</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>144,67,170,67</points>
<connection>
<GID>655</GID>
<name>N_in0</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>762</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,7.5,144.5,65.5</points>
<intersection>7.5 1</intersection>
<intersection>65.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,7.5,144.5,7.5</points>
<connection>
<GID>415</GID>
<name>OUT_5</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>144.5,65.5,170,65.5</points>
<connection>
<GID>654</GID>
<name>N_in0</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>763</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,6.5,145,64.5</points>
<intersection>6.5 1</intersection>
<intersection>64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,6.5,145,6.5</points>
<connection>
<GID>415</GID>
<name>OUT_4</name></connection>
<intersection>145 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>145,64.5,170,64.5</points>
<connection>
<GID>638</GID>
<name>N_in0</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>764</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,0,258,67.5</points>
<intersection>0 2</intersection>
<intersection>67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,67.5,267.5,67.5</points>
<connection>
<GID>664</GID>
<name>N_in0</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>145,0,258,0</points>
<intersection>145 3</intersection>
<intersection>258 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>145,0,145,5.5</points>
<intersection>0 2</intersection>
<intersection>5.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>143,5.5,145,5.5</points>
<connection>
<GID>415</GID>
<name>OUT_3</name></connection>
<intersection>145 3</intersection></hsegment></shape></wire>
<wire>
<ID>765</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,-1,259.5,66</points>
<intersection>-1 1</intersection>
<intersection>66 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-1,259.5,-1</points>
<intersection>144.5 3</intersection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,66,267.5,66</points>
<connection>
<GID>663</GID>
<name>N_in0</name></connection>
<intersection>259.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>144.5,-1,144.5,4.5</points>
<intersection>-1 1</intersection>
<intersection>4.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>143,4.5,144.5,4.5</points>
<connection>
<GID>415</GID>
<name>OUT_2</name></connection>
<intersection>144.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>766</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-2,261,64.5</points>
<intersection>-2 1</intersection>
<intersection>64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-2,261,-2</points>
<intersection>144 3</intersection>
<intersection>261 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>261,64.5,267.5,64.5</points>
<connection>
<GID>662</GID>
<name>N_in0</name></connection>
<intersection>261 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>144,-2,144,3.5</points>
<intersection>-2 1</intersection>
<intersection>3.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>143,3.5,144,3.5</points>
<connection>
<GID>415</GID>
<name>OUT_1</name></connection>
<intersection>144 3</intersection></hsegment></shape></wire>
<wire>
<ID>767</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263,-3.5,263,63.5</points>
<intersection>-3.5 1</intersection>
<intersection>63.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143.5,-3.5,263,-3.5</points>
<intersection>143.5 3</intersection>
<intersection>263 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>263,63.5,267.5,63.5</points>
<connection>
<GID>661</GID>
<name>N_in0</name></connection>
<intersection>263 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>143.5,-3.5,143.5,2.5</points>
<intersection>-3.5 1</intersection>
<intersection>2.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>143,2.5,143.5,2.5</points>
<connection>
<GID>415</GID>
<name>OUT_0</name></connection>
<intersection>143.5 3</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>243.451,157.487,984.177,-228.707</PageViewport>
<gate>
<ID>389</ID>
<type>AI_XOR2</type>
<position>334,-63</position>
<input>
<ID>IN_0</ID>530 </input>
<input>
<ID>IN_1</ID>543 </input>
<output>
<ID>OUT</ID>532 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>390</ID>
<type>AI_XOR2</type>
<position>338,-63</position>
<input>
<ID>IN_0</ID>530 </input>
<input>
<ID>IN_1</ID>542 </input>
<output>
<ID>OUT</ID>531 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>391</ID>
<type>AE_FULLADDER_4BIT</type>
<position>327,-74</position>
<input>
<ID>IN_1</ID>530 </input>
<input>
<ID>IN_3</ID>530 </input>
<input>
<ID>IN_B_0</ID>531 </input>
<input>
<ID>IN_B_1</ID>532 </input>
<input>
<ID>IN_B_2</ID>533 </input>
<input>
<ID>IN_B_3</ID>534 </input>
<output>
<ID>OUT_0</ID>541 </output>
<output>
<ID>OUT_1</ID>540 </output>
<output>
<ID>OUT_2</ID>539 </output>
<output>
<ID>OUT_3</ID>538 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>392</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>333.5,-83.5</position>
<input>
<ID>IN_0</ID>541 </input>
<input>
<ID>IN_1</ID>540 </input>
<input>
<ID>IN_2</ID>539 </input>
<input>
<ID>IN_3</ID>538 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>393</ID>
<type>GA_LED</type>
<position>324,-82.5</position>
<input>
<ID>N_in0</ID>535 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>394</ID>
<type>GA_LED</type>
<position>322,-82.5</position>
<input>
<ID>N_in0</ID>536 </input>
<input>
<ID>N_in1</ID>535 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>395</ID>
<type>GA_LED</type>
<position>320,-82.5</position>
<input>
<ID>N_in0</ID>537 </input>
<input>
<ID>N_in1</ID>536 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>396</ID>
<type>GA_LED</type>
<position>318,-82.5</position>
<input>
<ID>N_in0</ID>530 </input>
<input>
<ID>N_in1</ID>537 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>397</ID>
<type>AE_SMALL_INVERTER</type>
<position>314.5,-54.5</position>
<input>
<ID>IN_0</ID>352 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>398</ID>
<type>AI_XOR2</type>
<position>326,-37</position>
<input>
<ID>IN_0</ID>550 </input>
<input>
<ID>IN_1</ID>547 </input>
<output>
<ID>OUT</ID>546 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>399</ID>
<type>EE_VDD</type>
<position>325,-33</position>
<output>
<ID>OUT_0</ID>547 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>400</ID>
<type>AE_OR2</type>
<position>349,-49.5</position>
<input>
<ID>IN_0</ID>549 </input>
<input>
<ID>IN_1</ID>357 </input>
<output>
<ID>OUT</ID>358 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>401</ID>
<type>DD_KEYPAD_HEX</type>
<position>470.5,5.5</position>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>402</ID>
<type>DD_KEYPAD_HEX</type>
<position>470.5,17.5</position>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>403</ID>
<type>AA_AND2</type>
<position>531,30.5</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>372 </input>
<output>
<ID>OUT</ID>374 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_FULLADDER_4BIT</type>
<position>76,-35.5</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_3</ID>260 </input>
<input>
<ID>IN_B_0</ID>259 </input>
<input>
<ID>IN_B_1</ID>217 </input>
<input>
<ID>IN_B_2</ID>124 </input>
<input>
<ID>IN_B_3</ID>97 </input>
<output>
<ID>OUT_0</ID>76 </output>
<output>
<ID>OUT_1</ID>27 </output>
<output>
<ID>OUT_2</ID>26 </output>
<output>
<ID>OUT_3</ID>75 </output>
<input>
<ID>carry_in</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>404</ID>
<type>AA_AND2</type>
<position>531,19.5</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>371 </input>
<output>
<ID>OUT</ID>380 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>405</ID>
<type>AA_AND2</type>
<position>531,14</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>370 </input>
<output>
<ID>OUT</ID>402 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_AND2</type>
<position>531,9.5</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>369 </input>
<output>
<ID>OUT</ID>408 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>DD_KEYPAD_HEX</type>
<position>52,-33.5</position>
<output>
<ID>OUT_0</ID>273 </output>
<output>
<ID>OUT_1</ID>272 </output>
<output>
<ID>OUT_2</ID>271 </output>
<output>
<ID>OUT_3</ID>270 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>407</ID>
<type>AA_AND2</type>
<position>531,0</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>368 </input>
<output>
<ID>OUT</ID>410 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>63,-7</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_AND2</type>
<position>531,-4</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>351 </input>
<output>
<ID>OUT</ID>411 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>DD_KEYPAD_HEX</type>
<position>25.5,-47</position>
<output>
<ID>OUT_0</ID>106 </output>
<output>
<ID>OUT_1</ID>111 </output>
<output>
<ID>OUT_2</ID>118 </output>
<output>
<ID>OUT_3</ID>119 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_AND2</type>
<position>531,-8</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>350 </input>
<output>
<ID>OUT</ID>412 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>410</ID>
<type>AA_AND2</type>
<position>531,-12</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>314 </input>
<output>
<ID>OUT</ID>414 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>411</ID>
<type>AE_FULLADDER_4BIT</type>
<position>549.5,25.5</position>
<input>
<ID>IN_0</ID>442 </input>
<input>
<ID>IN_1</ID>441 </input>
<input>
<ID>IN_2</ID>440 </input>
<input>
<ID>IN_3</ID>425 </input>
<input>
<ID>IN_B_0</ID>374 </input>
<input>
<ID>IN_B_1</ID>380 </input>
<input>
<ID>IN_B_2</ID>402 </input>
<input>
<ID>IN_B_3</ID>408 </input>
<output>
<ID>OUT_0</ID>552 </output>
<output>
<ID>OUT_1</ID>551 </output>
<output>
<ID>OUT_2</ID>548 </output>
<output>
<ID>OUT_3</ID>522 </output>
<output>
<ID>carry_out</ID>553 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_FULLADDER_4BIT</type>
<position>84,-39</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>111 </input>
<input>
<ID>IN_2</ID>118 </input>
<input>
<ID>IN_3</ID>119 </input>
<input>
<ID>IN_B_0</ID>76 </input>
<input>
<ID>IN_B_1</ID>27 </input>
<input>
<ID>IN_B_2</ID>26 </input>
<input>
<ID>IN_B_3</ID>75 </input>
<output>
<ID>OUT_0</ID>59 </output>
<output>
<ID>OUT_1</ID>61 </output>
<output>
<ID>OUT_2</ID>60 </output>
<output>
<ID>OUT_3</ID>62 </output>
<output>
<ID>carry_out</ID>131 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>412</ID>
<type>AE_FULLADDER_4BIT</type>
<position>549.5,3.5</position>
<input>
<ID>IN_0</ID>424 </input>
<input>
<ID>IN_1</ID>423 </input>
<input>
<ID>IN_2</ID>422 </input>
<input>
<ID>IN_3</ID>417 </input>
<input>
<ID>IN_B_0</ID>410 </input>
<input>
<ID>IN_B_1</ID>411 </input>
<input>
<ID>IN_B_2</ID>412 </input>
<input>
<ID>IN_B_3</ID>414 </input>
<output>
<ID>OUT_0</ID>521 </output>
<output>
<ID>OUT_1</ID>519 </output>
<output>
<ID>OUT_2</ID>516 </output>
<output>
<ID>OUT_3</ID>481 </output>
<input>
<ID>carry_in</ID>553 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>413</ID>
<type>EE_VDD</type>
<position>533.5,-13.5</position>
<output>
<ID>OUT_0</ID>477 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_FULLADDER_4BIT</type>
<position>143,-26</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>210 </input>
<input>
<ID>IN_2</ID>209 </input>
<input>
<ID>IN_3</ID>216 </input>
<input>
<ID>IN_B_0</ID>59 </input>
<input>
<ID>IN_B_1</ID>61 </input>
<input>
<ID>IN_B_2</ID>60 </input>
<input>
<ID>IN_B_3</ID>62 </input>
<output>
<ID>OUT_0</ID>149 </output>
<output>
<ID>OUT_1</ID>148 </output>
<output>
<ID>OUT_2</ID>147 </output>
<output>
<ID>OUT_3</ID>146 </output>
<input>
<ID>carry_in</ID>260 </input>
<output>
<ID>carry_out</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>37</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>117,-42.5</position>
<output>
<ID>A_less_B</ID>151 </output>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_B_0</ID>59 </input>
<input>
<ID>IN_B_1</ID>61 </input>
<input>
<ID>IN_B_2</ID>60 </input>
<input>
<ID>IN_B_3</ID>62 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>39</ID>
<type>EE_VDD</type>
<position>107,-47.5</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>EE_VDD</type>
<position>107.5,-44.5</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>41</ID>
<type>AE_FULLADDER_4BIT</type>
<position>76,-75.5</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_3</ID>260 </input>
<input>
<ID>IN_B_0</ID>274 </input>
<input>
<ID>IN_B_1</ID>278 </input>
<input>
<ID>IN_B_2</ID>280 </input>
<input>
<ID>IN_B_3</ID>281 </input>
<output>
<ID>OUT_0</ID>263 </output>
<output>
<ID>OUT_1</ID>264 </output>
<output>
<ID>OUT_2</ID>262 </output>
<output>
<ID>OUT_3</ID>266 </output>
<input>
<ID>carry_in</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>53,-6.5</position>
<gparam>LABEL_TEXT is minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>61,-7</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>74.5,-6</position>
<gparam>LABEL_TEXT pressd minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AI_XOR2</type>
<position>-101.5,-25.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>421 </input>
<output>
<ID>OUT</ID>431 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AI_XOR2</type>
<position>62,-12</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>260 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AI_XOR2</type>
<position>-101.5,-29.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>420 </input>
<output>
<ID>OUT</ID>432 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_FULLADDER_4BIT</type>
<position>143,-63</position>
<input>
<ID>IN_0</ID>267 </input>
<input>
<ID>IN_1</ID>268 </input>
<input>
<ID>IN_2</ID>269 </input>
<input>
<ID>IN_3</ID>265 </input>
<input>
<ID>IN_B_0</ID>112 </input>
<input>
<ID>IN_B_1</ID>114 </input>
<input>
<ID>IN_B_2</ID>113 </input>
<input>
<ID>IN_B_3</ID>115 </input>
<output>
<ID>OUT_0</ID>157 </output>
<output>
<ID>OUT_1</ID>158 </output>
<output>
<ID>OUT_2</ID>159 </output>
<output>
<ID>OUT_3</ID>161 </output>
<input>
<ID>carry_in</ID>164 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>55</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>120.5,-78</position>
<output>
<ID>A_less_B</ID>162 </output>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_3</ID>116 </input>
<input>
<ID>IN_B_0</ID>112 </input>
<input>
<ID>IN_B_1</ID>114 </input>
<input>
<ID>IN_B_2</ID>113 </input>
<input>
<ID>IN_B_3</ID>115 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>61</ID>
<type>EE_VDD</type>
<position>115.5,-83</position>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>DD_KEYPAD_HEX</type>
<position>212,-38.5</position>
<output>
<ID>OUT_0</ID>35 </output>
<output>
<ID>OUT_1</ID>36 </output>
<output>
<ID>OUT_2</ID>37 </output>
<output>
<ID>OUT_3</ID>38 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>63</ID>
<type>GA_LED</type>
<position>166.5,-74.5</position>
<input>
<ID>N_in2</ID>121 </input>
<input>
<ID>N_in3</ID>207 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>DD_KEYPAD_HEX</type>
<position>185.5,-50.5</position>
<output>
<ID>OUT_0</ID>49 </output>
<output>
<ID>OUT_1</ID>48 </output>
<output>
<ID>OUT_2</ID>47 </output>
<output>
<ID>OUT_3</ID>46 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_FULLADDER_4BIT</type>
<position>240,-44</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>48 </input>
<input>
<ID>IN_2</ID>47 </input>
<input>
<ID>IN_3</ID>46 </input>
<input>
<ID>IN_B_0</ID>35 </input>
<input>
<ID>IN_B_1</ID>36 </input>
<input>
<ID>IN_B_2</ID>37 </input>
<input>
<ID>IN_B_3</ID>38 </input>
<output>
<ID>OUT_0</ID>39 </output>
<output>
<ID>OUT_1</ID>41 </output>
<output>
<ID>OUT_2</ID>40 </output>
<output>
<ID>OUT_3</ID>42 </output>
<output>
<ID>carry_out</ID>153 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>67</ID>
<type>AE_FULLADDER_4BIT</type>
<position>289,-31</position>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>50 </input>
<input>
<ID>IN_B_0</ID>39 </input>
<input>
<ID>IN_B_1</ID>41 </input>
<input>
<ID>IN_B_2</ID>40 </input>
<input>
<ID>IN_B_3</ID>42 </input>
<output>
<ID>OUT_0</ID>172 </output>
<output>
<ID>OUT_1</ID>171 </output>
<output>
<ID>OUT_2</ID>165 </output>
<output>
<ID>OUT_3</ID>156 </output>
<output>
<ID>carry_out</ID>201 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>70</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>165,-26.5</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>148 </input>
<input>
<ID>IN_2</ID>147 </input>
<input>
<ID>IN_3</ID>146 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_OR2</type>
<position>122.5,-47.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>208 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>166.5,-63.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>158 </input>
<input>
<ID>IN_2</ID>159 </input>
<input>
<ID>IN_3</ID>161 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_OR2</type>
<position>126,-89.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>296 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>277,-47.5</position>
<output>
<ID>A_less_B</ID>173 </output>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_3</ID>43 </input>
<input>
<ID>IN_B_0</ID>39 </input>
<input>
<ID>IN_B_1</ID>41 </input>
<input>
<ID>IN_B_2</ID>40 </input>
<input>
<ID>IN_B_3</ID>42 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>76</ID>
<type>EE_VDD</type>
<position>267,-52.5</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>77</ID>
<type>EE_VDD</type>
<position>267.5,-49.5</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>78</ID>
<type>AI_XOR2</type>
<position>112,-80</position>
<input>
<ID>IN_0</ID>166 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AI_XOR2</type>
<position>-101.5,-33.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>419 </input>
<output>
<ID>OUT</ID>433 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>EE_VDD</type>
<position>108,-79</position>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>166.5,-76.5</position>
<input>
<ID>N_in2</ID>123 </input>
<input>
<ID>N_in3</ID>121 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AI_XOR2</type>
<position>-101.5,-37.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>418 </input>
<output>
<ID>OUT</ID>434 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>DD_KEYPAD_HEX</type>
<position>212.5,-75</position>
<output>
<ID>OUT_0</ID>51 </output>
<output>
<ID>OUT_1</ID>53 </output>
<output>
<ID>OUT_2</ID>57 </output>
<output>
<ID>OUT_3</ID>58 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>DD_KEYPAD_HEX</type>
<position>188,-87</position>
<output>
<ID>OUT_0</ID>137 </output>
<output>
<ID>OUT_1</ID>127 </output>
<output>
<ID>OUT_2</ID>126 </output>
<output>
<ID>OUT_3</ID>125 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>85</ID>
<type>AE_FULLADDER_4BIT</type>
<position>240,-79.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>127 </input>
<input>
<ID>IN_2</ID>126 </input>
<input>
<ID>IN_3</ID>125 </input>
<input>
<ID>IN_B_0</ID>51 </input>
<input>
<ID>IN_B_1</ID>53 </input>
<input>
<ID>IN_B_2</ID>57 </input>
<input>
<ID>IN_B_3</ID>58 </input>
<output>
<ID>OUT_0</ID>74 </output>
<output>
<ID>OUT_1</ID>101 </output>
<output>
<ID>OUT_2</ID>98 </output>
<output>
<ID>OUT_3</ID>102 </output>
<input>
<ID>carry_in</ID>153 </input>
<output>
<ID>carry_out</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>86</ID>
<type>AE_FULLADDER_4BIT</type>
<position>291.5,-68</position>
<input>
<ID>IN_1</ID>150 </input>
<input>
<ID>IN_2</ID>150 </input>
<input>
<ID>IN_B_0</ID>74 </input>
<input>
<ID>IN_B_1</ID>101 </input>
<input>
<ID>IN_B_2</ID>98 </input>
<input>
<ID>IN_B_3</ID>102 </input>
<output>
<ID>OUT_0</ID>180 </output>
<output>
<ID>OUT_1</ID>182 </output>
<output>
<ID>OUT_2</ID>183 </output>
<output>
<ID>OUT_3</ID>184 </output>
<input>
<ID>carry_in</ID>201 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>92</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>280.5,-83</position>
<output>
<ID>A_less_B</ID>185 </output>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_3</ID>103 </input>
<input>
<ID>IN_B_0</ID>74 </input>
<input>
<ID>IN_B_1</ID>101 </input>
<input>
<ID>IN_B_2</ID>98 </input>
<input>
<ID>IN_B_3</ID>102 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>93</ID>
<type>EE_VDD</type>
<position>275.5,-88</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>114</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>302,-31</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>171 </input>
<input>
<ID>IN_2</ID>165 </input>
<input>
<ID>IN_3</ID>156 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 8</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_OR2</type>
<position>283.5,-53</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>303.5,-68.5</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>182 </input>
<input>
<ID>IN_2</ID>183 </input>
<input>
<ID>IN_3</ID>184 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_OR2</type>
<position>286,-94.5</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>200 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>AI_XOR2</type>
<position>272,-85</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>201 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>EE_VDD</type>
<position>268,-84</position>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>129</ID>
<type>GA_LED</type>
<position>166.5,-78.5</position>
<input>
<ID>N_in0</ID>163 </input>
<input>
<ID>N_in2</ID>163 </input>
<input>
<ID>N_in3</ID>123 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>FF_GND</type>
<position>-37,-29.5</position>
<output>
<ID>OUT_0</ID>403 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>173</ID>
<type>FF_GND</type>
<position>-37,-41.5</position>
<output>
<ID>OUT_0</ID>404 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>174</ID>
<type>GA_LED</type>
<position>166.5,-80.5</position>
<input>
<ID>N_in3</ID>163 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>FF_GND</type>
<position>-36.5,-65.5</position>
<output>
<ID>OUT_0</ID>406 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_AND2</type>
<position>82,-9.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>AI_XOR2</type>
<position>134.5,-27</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>219 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>190</ID>
<type>AI_XOR2</type>
<position>134.5,-31</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>AI_XOR2</type>
<position>134.5,-35</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>AI_XOR2</type>
<position>134.5,-39</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>221 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>193</ID>
<type>FF_GND</type>
<position>-36.5,-77.5</position>
<output>
<ID>OUT_0</ID>407 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>195</ID>
<type>AI_XOR2</type>
<position>66,-24</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>273 </input>
<output>
<ID>OUT</ID>259 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>198</ID>
<type>AI_XOR2</type>
<position>66,-28</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AI_XOR2</type>
<position>66,-32</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>271 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>AI_XOR2</type>
<position>66,-36</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>270 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>FF_GND</type>
<position>130.5,-28</position>
<output>
<ID>OUT_0</ID>219 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>202</ID>
<type>FF_GND</type>
<position>130.5,-40</position>
<output>
<ID>OUT_0</ID>221 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>203</ID>
<type>FF_GND</type>
<position>131,-64</position>
<output>
<ID>OUT_0</ID>252 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>204</ID>
<type>FF_GND</type>
<position>131,-76</position>
<output>
<ID>OUT_0</ID>253 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>206</ID>
<type>AI_XOR2</type>
<position>65,-65</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>291 </input>
<output>
<ID>OUT</ID>274 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>AI_XOR2</type>
<position>65,-69</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>290 </input>
<output>
<ID>OUT</ID>278 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>208</ID>
<type>AI_XOR2</type>
<position>65,-73</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>289 </input>
<output>
<ID>OUT</ID>280 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>209</ID>
<type>AI_XOR2</type>
<position>65,-77</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>288 </input>
<output>
<ID>OUT</ID>281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>AI_XOR2</type>
<position>135,-63</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>AI_XOR2</type>
<position>135,-67</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>AI_XOR2</type>
<position>135,-71</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>269 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>AI_XOR2</type>
<position>135,-75</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>253 </input>
<output>
<ID>OUT</ID>265 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>DD_KEYPAD_HEX</type>
<position>50.5,-74.5</position>
<output>
<ID>OUT_0</ID>291 </output>
<output>
<ID>OUT_1</ID>290 </output>
<output>
<ID>OUT_2</ID>289 </output>
<output>
<ID>OUT_3</ID>288 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>215</ID>
<type>AI_XOR2</type>
<position>-102.5,-66.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>429 </input>
<output>
<ID>OUT</ID>435 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>DD_KEYPAD_HEX</type>
<position>26,-88</position>
<output>
<ID>OUT_0</ID>105 </output>
<output>
<ID>OUT_1</ID>104 </output>
<output>
<ID>OUT_2</ID>96 </output>
<output>
<ID>OUT_3</ID>95 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>217</ID>
<type>AE_FULLADDER_4BIT</type>
<position>84,-79</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>104 </input>
<input>
<ID>IN_2</ID>96 </input>
<input>
<ID>IN_3</ID>95 </input>
<input>
<ID>IN_B_0</ID>263 </input>
<input>
<ID>IN_B_1</ID>264 </input>
<input>
<ID>IN_B_2</ID>262 </input>
<input>
<ID>IN_B_3</ID>266 </input>
<output>
<ID>OUT_0</ID>112 </output>
<output>
<ID>OUT_1</ID>114 </output>
<output>
<ID>OUT_2</ID>113 </output>
<output>
<ID>OUT_3</ID>115 </output>
<input>
<ID>carry_in</ID>131 </input>
<output>
<ID>carry_out</ID>296 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>218</ID>
<type>AI_XOR2</type>
<position>381.5,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>325 </input>
<output>
<ID>OUT</ID>279 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>AI_XOR2</type>
<position>385.5,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>326 </input>
<output>
<ID>OUT</ID>277 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>AI_XOR2</type>
<position>389.5,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>327 </input>
<output>
<ID>OUT</ID>276 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>AI_XOR2</type>
<position>393.5,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>328 </input>
<output>
<ID>OUT</ID>275 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>30,-28</position>
<gparam>LABEL_TEXT /</gparam>
<gparam>TEXT_HEIGHT 12</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>DD_KEYPAD_HEX</type>
<position>490,21.5</position>
<output>
<ID>OUT_0</ID>558 </output>
<output>
<ID>OUT_1</ID>557 </output>
<output>
<ID>OUT_2</ID>556 </output>
<output>
<ID>OUT_3</ID>555 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>224</ID>
<type>AI_XOR2</type>
<position>-102.5,-70.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>428 </input>
<output>
<ID>OUT</ID>436 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>AI_XOR2</type>
<position>-102.5,-74.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>427 </input>
<output>
<ID>OUT</ID>437 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>226</ID>
<type>AI_XOR2</type>
<position>-102.5,-78.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>426 </input>
<output>
<ID>OUT</ID>438 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>DD_KEYPAD_HEX</type>
<position>-115.5,-35</position>
<output>
<ID>OUT_0</ID>421 </output>
<output>
<ID>OUT_1</ID>420 </output>
<output>
<ID>OUT_2</ID>419 </output>
<output>
<ID>OUT_3</ID>418 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 4</lparam></gate>
<gate>
<ID>228</ID>
<type>AE_FULLADDER_4BIT</type>
<position>379.5,-15.5</position>
<input>
<ID>IN_1</ID>292 </input>
<input>
<ID>IN_3</ID>292 </input>
<input>
<ID>IN_B_0</ID>275 </input>
<input>
<ID>IN_B_1</ID>276 </input>
<input>
<ID>IN_B_2</ID>277 </input>
<input>
<ID>IN_B_3</ID>279 </input>
<output>
<ID>OUT_0</ID>297 </output>
<output>
<ID>OUT_1</ID>299 </output>
<output>
<ID>OUT_2</ID>295 </output>
<output>
<ID>OUT_3</ID>298 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>229</ID>
<type>AI_XOR2</type>
<position>-32.5,-64.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>406 </input>
<output>
<ID>OUT</ID>415 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_TOGGLE</type>
<position>-104.5,-8.5</position>
<output>
<ID>OUT_0</ID>284 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>231</ID>
<type>AI_XOR2</type>
<position>-32.5,-68.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>405 </input>
<output>
<ID>OUT</ID>416 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>232</ID>
<type>DD_KEYPAD_HEX</type>
<position>-142.5,-48.5</position>
<output>
<ID>OUT_0</ID>341 </output>
<output>
<ID>OUT_1</ID>344 </output>
<output>
<ID>OUT_2</ID>376 </output>
<output>
<ID>OUT_3</ID>377 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>233</ID>
<type>AI_XOR2</type>
<position>-32.5,-72.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>405 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>234</ID>
<type>AI_XOR2</type>
<position>-32.5,-76.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>407 </input>
<output>
<ID>OUT</ID>413 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>235</ID>
<type>DD_KEYPAD_HEX</type>
<position>-117,-76</position>
<output>
<ID>OUT_0</ID>429 </output>
<output>
<ID>OUT_1</ID>428 </output>
<output>
<ID>OUT_2</ID>427 </output>
<output>
<ID>OUT_3</ID>426 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>236</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-83.5,-40.5</position>
<input>
<ID>IN_0</ID>341 </input>
<input>
<ID>IN_1</ID>344 </input>
<input>
<ID>IN_2</ID>376 </input>
<input>
<ID>IN_3</ID>377 </input>
<input>
<ID>IN_B_0</ID>431 </input>
<input>
<ID>IN_B_1</ID>432 </input>
<input>
<ID>IN_B_2</ID>433 </input>
<input>
<ID>IN_B_3</ID>434 </input>
<output>
<ID>OUT_0</ID>287 </output>
<output>
<ID>OUT_1</ID>294 </output>
<output>
<ID>OUT_2</ID>293 </output>
<output>
<ID>OUT_3</ID>300 </output>
<input>
<ID>carry_in</ID>409 </input>
<output>
<ID>carry_out</ID>381 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>238</ID>
<type>DD_KEYPAD_HEX</type>
<position>-141.5,-89.5</position>
<output>
<ID>OUT_0</ID>320 </output>
<output>
<ID>OUT_1</ID>319 </output>
<output>
<ID>OUT_2</ID>309 </output>
<output>
<ID>OUT_3</ID>308 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>240</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-83.5,-80.5</position>
<input>
<ID>IN_0</ID>320 </input>
<input>
<ID>IN_1</ID>319 </input>
<input>
<ID>IN_2</ID>309 </input>
<input>
<ID>IN_3</ID>308 </input>
<input>
<ID>IN_B_0</ID>435 </input>
<input>
<ID>IN_B_1</ID>436 </input>
<input>
<ID>IN_B_2</ID>437 </input>
<input>
<ID>IN_B_3</ID>438 </input>
<output>
<ID>OUT_0</ID>354 </output>
<output>
<ID>OUT_1</ID>356 </output>
<output>
<ID>OUT_2</ID>355 </output>
<output>
<ID>OUT_3</ID>363 </output>
<input>
<ID>carry_in</ID>381 </input>
<output>
<ID>carry_out</ID>430 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_FULLADDER_4BIT</type>
<position>370.5,-29</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>331 </input>
<input>
<ID>IN_2</ID>330 </input>
<input>
<ID>IN_3</ID>329 </input>
<input>
<ID>IN_B_0</ID>297 </input>
<input>
<ID>IN_B_1</ID>299 </input>
<input>
<ID>IN_B_2</ID>295 </input>
<input>
<ID>IN_B_3</ID>298 </input>
<output>
<ID>OUT_0</ID>339 </output>
<output>
<ID>OUT_1</ID>338 </output>
<output>
<ID>OUT_2</ID>337 </output>
<output>
<ID>OUT_3</ID>340 </output>
<output>
<ID>carry_out</ID>357 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>242</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-24.5,-27.5</position>
<input>
<ID>IN_0</ID>400 </input>
<input>
<ID>IN_1</ID>399 </input>
<input>
<ID>IN_2</ID>398 </input>
<input>
<ID>IN_3</ID>401 </input>
<input>
<ID>IN_B_0</ID>287 </input>
<input>
<ID>IN_B_1</ID>294 </input>
<input>
<ID>IN_B_2</ID>293 </input>
<input>
<ID>IN_B_3</ID>300 </input>
<output>
<ID>OUT_0</ID>385 </output>
<output>
<ID>OUT_1</ID>384 </output>
<output>
<ID>OUT_2</ID>383 </output>
<output>
<ID>OUT_3</ID>382 </output>
<input>
<ID>carry_in</ID>409 </input>
<output>
<ID>carry_out</ID>393 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>244</ID>
<type>DD_KEYPAD_HEX</type>
<position>344,24.5</position>
<output>
<ID>OUT_0</ID>336 </output>
<output>
<ID>OUT_1</ID>335 </output>
<output>
<ID>OUT_2</ID>334 </output>
<output>
<ID>OUT_3</ID>333 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>245</ID>
<type>DD_KEYPAD_HEX</type>
<position>355.5,24.5</position>
<output>
<ID>OUT_0</ID>332 </output>
<output>
<ID>OUT_1</ID>331 </output>
<output>
<ID>OUT_2</ID>330 </output>
<output>
<ID>OUT_3</ID>329 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>246</ID>
<type>DD_KEYPAD_HEX</type>
<position>376.5,24.5</position>
<output>
<ID>OUT_0</ID>324 </output>
<output>
<ID>OUT_1</ID>323 </output>
<output>
<ID>OUT_2</ID>322 </output>
<output>
<ID>OUT_3</ID>321 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>248</ID>
<type>DD_KEYPAD_HEX</type>
<position>391,24</position>
<output>
<ID>OUT_0</ID>328 </output>
<output>
<ID>OUT_1</ID>327 </output>
<output>
<ID>OUT_2</ID>326 </output>
<output>
<ID>OUT_3</ID>325 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_LABEL</type>
<position>-137.5,-29.5</position>
<gparam>LABEL_TEXT /</gparam>
<gparam>TEXT_HEIGHT 12</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>GA_LED</type>
<position>276,6.5</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>-50.5,-44</position>
<output>
<ID>A_less_B</ID>386 </output>
<input>
<ID>IN_0</ID>302 </input>
<input>
<ID>IN_3</ID>301 </input>
<input>
<ID>IN_B_0</ID>287 </input>
<input>
<ID>IN_B_1</ID>294 </input>
<input>
<ID>IN_B_2</ID>293 </input>
<input>
<ID>IN_B_3</ID>300 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_TOGGLE</type>
<position>305.5,14</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>254</ID>
<type>EE_VDD</type>
<position>-60.5,-49</position>
<output>
<ID>OUT_0</ID>301 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>257</ID>
<type>CC_PULSE</type>
<position>355,38.5</position>
<output>
<ID>OUT_0</ID>306 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>EE_VDD</type>
<position>-60,-46</position>
<output>
<ID>OUT_0</ID>302 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>259</ID>
<type>BE_JKFF_LOW</type>
<position>360,38.5</position>
<input>
<ID>J</ID>306 </input>
<input>
<ID>K</ID>306 </input>
<output>
<ID>Q</ID>305 </output>
<input>
<ID>clock</ID>306 </input>
<output>
<ID>nQ</ID>292 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>260</ID>
<type>DD_KEYPAD_HEX</type>
<position>489.5,5</position>
<output>
<ID>OUT_0</ID>562 </output>
<output>
<ID>OUT_1</ID>561 </output>
<output>
<ID>OUT_2</ID>560 </output>
<output>
<ID>OUT_3</ID>559 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>261</ID>
<type>GA_LED</type>
<position>366.5,24.5</position>
<input>
<ID>N_in1</ID>307 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>-114.5,-8</position>
<gparam>LABEL_TEXT is minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>264</ID>
<type>GA_LED</type>
<position>366.5,22.5</position>
<input>
<ID>N_in2</ID>305 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>265</ID>
<type>AA_TOGGLE</type>
<position>-106.5,-8.5</position>
<output>
<ID>OUT_0</ID>283 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>266</ID>
<type>GA_LED</type>
<position>366.5,26.5</position>
<input>
<ID>N_in1</ID>305 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>AA_LABEL</type>
<position>-93,-7.5</position>
<gparam>LABEL_TEXT pressd minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>268</ID>
<type>GA_LED</type>
<position>368.5,24.5</position>
<input>
<ID>N_in1</ID>307 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>271</ID>
<type>AI_XOR2</type>
<position>-105.5,-13.5</position>
<input>
<ID>IN_0</ID>284 </input>
<input>
<ID>IN_1</ID>283 </input>
<output>
<ID>OUT</ID>409 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>272</ID>
<type>GA_LED</type>
<position>364.5,24.5</position>
<input>
<ID>N_in1</ID>307 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>273</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-24.5,-64.5</position>
<input>
<ID>IN_0</ID>415 </input>
<input>
<ID>IN_1</ID>416 </input>
<input>
<ID>IN_3</ID>413 </input>
<input>
<ID>IN_B_0</ID>354 </input>
<input>
<ID>IN_B_1</ID>356 </input>
<input>
<ID>IN_B_2</ID>355 </input>
<input>
<ID>IN_B_3</ID>363 </input>
<output>
<ID>OUT_0</ID>387 </output>
<output>
<ID>OUT_1</ID>388 </output>
<output>
<ID>OUT_2</ID>389 </output>
<output>
<ID>OUT_3</ID>390 </output>
<input>
<ID>carry_in</ID>393 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>274</ID>
<type>AE_OR2</type>
<position>366.5,34.5</position>
<input>
<ID>IN_0</ID>305 </input>
<input>
<ID>IN_1</ID>292 </input>
<output>
<ID>OUT</ID>307 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>-47,-79.5</position>
<output>
<ID>A_less_B</ID>391 </output>
<input>
<ID>IN_0</ID>395 </input>
<input>
<ID>IN_3</ID>375 </input>
<input>
<ID>IN_B_0</ID>354 </input>
<input>
<ID>IN_B_1</ID>356 </input>
<input>
<ID>IN_B_2</ID>355 </input>
<input>
<ID>IN_B_3</ID>363 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_LABEL</type>
<position>409,4.5</position>
<gparam>LABEL_TEXT minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>277</ID>
<type>AI_XOR2</type>
<position>350,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>321 </input>
<output>
<ID>OUT</ID>313 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>AI_XOR2</type>
<position>354,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>312 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>AI_XOR2</type>
<position>358,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>323 </input>
<output>
<ID>OUT</ID>311 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>670</ID>
<type>BB_CLOCK</type>
<position>491.5,-23</position>
<output>
<ID>CLK</ID>303 </output>
<gparam>angle 0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>281</ID>
<type>AI_XOR2</type>
<position>362,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>324 </input>
<output>
<ID>OUT</ID>310 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>AE_FULLADDER_4BIT</type>
<position>348,-15.5</position>
<input>
<ID>IN_1</ID>292 </input>
<input>
<ID>IN_3</ID>292 </input>
<input>
<ID>IN_B_0</ID>310 </input>
<input>
<ID>IN_B_1</ID>311 </input>
<input>
<ID>IN_B_2</ID>312 </input>
<input>
<ID>IN_B_3</ID>313 </input>
<output>
<ID>OUT_0</ID>316 </output>
<output>
<ID>OUT_1</ID>318 </output>
<output>
<ID>OUT_2</ID>315 </output>
<output>
<ID>OUT_3</ID>317 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>672</ID>
<type>CC_PULSE</type>
<position>518,-20</position>
<output>
<ID>OUT_0</ID>261 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>283</ID>
<type>AE_FULLADDER_4BIT</type>
<position>339,-29</position>
<input>
<ID>IN_0</ID>336 </input>
<input>
<ID>IN_1</ID>335 </input>
<input>
<ID>IN_2</ID>334 </input>
<input>
<ID>IN_3</ID>333 </input>
<input>
<ID>IN_B_0</ID>316 </input>
<input>
<ID>IN_B_1</ID>318 </input>
<input>
<ID>IN_B_2</ID>315 </input>
<input>
<ID>IN_B_3</ID>317 </input>
<output>
<ID>OUT_0</ID>347 </output>
<output>
<ID>OUT_1</ID>346 </output>
<output>
<ID>OUT_2</ID>345 </output>
<output>
<ID>OUT_3</ID>348 </output>
<input>
<ID>carry_in</ID>357 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>673</ID>
<type>CC_PULSE</type>
<position>515,-34.5</position>
<output>
<ID>OUT_0</ID>554 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>284</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>359.5,-44.5</position>
<output>
<ID>A_less_B</ID>549 </output>
<input>
<ID>IN_0</ID>343 </input>
<input>
<ID>IN_3</ID>342 </input>
<input>
<ID>IN_B_0</ID>339 </input>
<input>
<ID>IN_B_1</ID>338 </input>
<input>
<ID>IN_B_2</ID>337 </input>
<input>
<ID>IN_B_3</ID>340 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>285</ID>
<type>EE_VDD</type>
<position>-52,-84.5</position>
<output>
<ID>OUT_0</ID>375 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>286</ID>
<type>EE_VDD</type>
<position>354.5,-39.5</position>
<output>
<ID>OUT_0</ID>342 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>287</ID>
<type>EE_VDD</type>
<position>357.5,-39.5</position>
<output>
<ID>OUT_0</ID>343 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>288</ID>
<type>AE_FULLADDER_4BIT</type>
<position>367,-53</position>
<input>
<ID>IN_1</ID>358 </input>
<input>
<ID>IN_2</ID>358 </input>
<input>
<ID>IN_B_0</ID>339 </input>
<input>
<ID>IN_B_1</ID>338 </input>
<input>
<ID>IN_B_2</ID>337 </input>
<input>
<ID>IN_B_3</ID>340 </input>
<output>
<ID>OUT_0</ID>367 </output>
<output>
<ID>OUT_1</ID>366 </output>
<output>
<ID>OUT_2</ID>365 </output>
<output>
<ID>OUT_3</ID>364 </output>
<output>
<ID>carry_out</ID>550 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>290</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>328,-44</position>
<output>
<ID>A_less_B</ID>352 </output>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_3</ID>349 </input>
<input>
<ID>IN_B_0</ID>347 </input>
<input>
<ID>IN_B_1</ID>346 </input>
<input>
<ID>IN_B_2</ID>345 </input>
<input>
<ID>IN_B_3</ID>348 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>295</ID>
<type>EE_VDD</type>
<position>323,-39</position>
<output>
<ID>OUT_0</ID>349 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>297</ID>
<type>AE_FULLADDER_4BIT</type>
<position>335.5,-53</position>
<input>
<ID>IN_1</ID>352 </input>
<input>
<ID>IN_2</ID>352 </input>
<input>
<ID>IN_B_0</ID>347 </input>
<input>
<ID>IN_B_1</ID>346 </input>
<input>
<ID>IN_B_2</ID>345 </input>
<input>
<ID>IN_B_3</ID>348 </input>
<output>
<ID>OUT_0</ID>542 </output>
<output>
<ID>OUT_1</ID>543 </output>
<output>
<ID>OUT_2</ID>544 </output>
<output>
<ID>OUT_3</ID>545 </output>
<input>
<ID>carry_in</ID>550 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>298</ID>
<type>AI_XOR2</type>
<position>359.5,-63</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>362 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>299</ID>
<type>AI_XOR2</type>
<position>363.5,-63</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>365 </input>
<output>
<ID>OUT</ID>361 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>300</ID>
<type>AI_XOR2</type>
<position>367.5,-63</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>360 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>301</ID>
<type>AI_XOR2</type>
<position>371.5,-63</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>367 </input>
<output>
<ID>OUT</ID>359 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>AE_FULLADDER_4BIT</type>
<position>360.5,-74</position>
<input>
<ID>IN_1</ID>353 </input>
<input>
<ID>IN_3</ID>353 </input>
<input>
<ID>IN_B_0</ID>359 </input>
<input>
<ID>IN_B_1</ID>360 </input>
<input>
<ID>IN_B_2</ID>361 </input>
<input>
<ID>IN_B_3</ID>362 </input>
<output>
<ID>OUT_0</ID>529 </output>
<output>
<ID>OUT_1</ID>528 </output>
<output>
<ID>OUT_2</ID>527 </output>
<output>
<ID>OUT_3</ID>526 </output>
<input>
<ID>carry_in</ID>358 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>304</ID>
<type>GA_LED</type>
<position>-1,-76</position>
<input>
<ID>N_in2</ID>378 </input>
<input>
<ID>N_in3</ID>396 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>305</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-2.5,-28</position>
<input>
<ID>IN_0</ID>385 </input>
<input>
<ID>IN_1</ID>384 </input>
<input>
<ID>IN_2</ID>383 </input>
<input>
<ID>IN_3</ID>382 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_OR2</type>
<position>-45,-49</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>439 </input>
<output>
<ID>OUT</ID>397 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>AE_SMALL_INVERTER</type>
<position>349,-56.5</position>
<input>
<ID>IN_0</ID>358 </input>
<output>
<ID>OUT_0</ID>353 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>308</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>367,-83.5</position>
<input>
<ID>IN_0</ID>529 </input>
<input>
<ID>IN_1</ID>528 </input>
<input>
<ID>IN_2</ID>527 </input>
<input>
<ID>IN_3</ID>526 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>309</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-1,-65</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>388 </input>
<input>
<ID>IN_2</ID>389 </input>
<input>
<ID>IN_3</ID>390 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 12</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>310</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>589,-37.5</position>
<input>
<ID>IN_0</ID>552 </input>
<input>
<ID>IN_1</ID>551 </input>
<input>
<ID>IN_2</ID>548 </input>
<input>
<ID>IN_3</ID>522 </input>
<input>
<ID>IN_4</ID>521 </input>
<input>
<ID>IN_5</ID>519 </input>
<input>
<ID>IN_6</ID>516 </input>
<input>
<ID>IN_7</ID>481 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>311</ID>
<type>AE_REGISTER8</type>
<position>534,-22</position>
<input>
<ID>IN_0</ID>552 </input>
<input>
<ID>IN_1</ID>551 </input>
<input>
<ID>IN_2</ID>548 </input>
<input>
<ID>IN_3</ID>522 </input>
<input>
<ID>IN_4</ID>521 </input>
<input>
<ID>IN_5</ID>519 </input>
<input>
<ID>IN_6</ID>516 </input>
<input>
<ID>IN_7</ID>481 </input>
<output>
<ID>OUT_0</ID>442 </output>
<output>
<ID>OUT_1</ID>441 </output>
<output>
<ID>OUT_2</ID>440 </output>
<output>
<ID>OUT_3</ID>425 </output>
<output>
<ID>OUT_4</ID>424 </output>
<output>
<ID>OUT_5</ID>423 </output>
<output>
<ID>OUT_6</ID>422 </output>
<output>
<ID>OUT_7</ID>417 </output>
<input>
<ID>clear</ID>554 </input>
<input>
<ID>clock</ID>303 </input>
<input>
<ID>load</ID>477 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>312</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>511,27</position>
<input>
<ID>IN_0</ID>555 </input>
<input>
<ID>IN_1</ID>556 </input>
<input>
<ID>IN_2</ID>557 </input>
<input>
<ID>IN_3</ID>558 </input>
<output>
<ID>carry_out</ID>373 </output>
<input>
<ID>clear</ID>554 </input>
<input>
<ID>clock</ID>303 </input>
<input>
<ID>load</ID>261 </input>
<input>
<ID>shift_enable</ID>769 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>313</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>510,10</position>
<input>
<ID>IN_0</ID>562 </input>
<input>
<ID>IN_1</ID>561 </input>
<input>
<ID>IN_2</ID>560 </input>
<input>
<ID>IN_3</ID>559 </input>
<output>
<ID>OUT_0</ID>372 </output>
<output>
<ID>OUT_1</ID>371 </output>
<output>
<ID>OUT_2</ID>370 </output>
<output>
<ID>OUT_3</ID>369 </output>
<output>
<ID>carry_out</ID>304 </output>
<input>
<ID>clear</ID>554 </input>
<input>
<ID>clock</ID>303 </input>
<input>
<ID>load</ID>261 </input>
<input>
<ID>shift_enable</ID>768 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>314</ID>
<type>AE_OR2</type>
<position>-42,-91</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>430 </input>
<output>
<ID>OUT</ID>443 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>315</ID>
<type>AI_XOR2</type>
<position>-55.5,-81.5</position>
<input>
<ID>IN_0</ID>394 </input>
<input>
<ID>IN_1</ID>393 </input>
<output>
<ID>OUT</ID>395 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>316</ID>
<type>EE_VDD</type>
<position>-59.5,-80.5</position>
<output>
<ID>OUT_0</ID>394 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>317</ID>
<type>GA_LED</type>
<position>-1,-78</position>
<input>
<ID>N_in2</ID>379 </input>
<input>
<ID>N_in3</ID>378 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>318</ID>
<type>GA_LED</type>
<position>-1,-80</position>
<input>
<ID>N_in0</ID>392 </input>
<input>
<ID>N_in2</ID>392 </input>
<input>
<ID>N_in3</ID>379 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>319</ID>
<type>GA_LED</type>
<position>-1,-82</position>
<input>
<ID>N_in3</ID>392 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>320</ID>
<type>AA_AND2</type>
<position>-85.5,-11</position>
<input>
<ID>IN_0</ID>283 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>396 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>321</ID>
<type>AI_XOR2</type>
<position>-33,-28.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>403 </input>
<output>
<ID>OUT</ID>400 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>322</ID>
<type>AI_XOR2</type>
<position>-33,-32.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>399 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>323</ID>
<type>AI_XOR2</type>
<position>-33,-36.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>398 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>324</ID>
<type>AI_XOR2</type>
<position>-33,-40.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>404 </input>
<output>
<ID>OUT</ID>401 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>325</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>510,-6</position>
<output>
<ID>OUT_0</ID>368 </output>
<output>
<ID>OUT_1</ID>351 </output>
<output>
<ID>OUT_2</ID>350 </output>
<output>
<ID>OUT_3</ID>314 </output>
<input>
<ID>carry_in</ID>304 </input>
<input>
<ID>clear</ID>554 </input>
<input>
<ID>clock</ID>303 </input>
<input>
<ID>load</ID>261 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>326</ID>
<type>AI_XOR2</type>
<position>-72.5,-54</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>381 </input>
<output>
<ID>OUT</ID>439 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>AI_XOR2</type>
<position>-36,-84.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>443 </input>
<output>
<ID>OUT</ID>405 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>330</ID>
<type>FF_GND</type>
<position>-198,-79.5</position>
<output>
<ID>OUT_0</ID>492 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>331</ID>
<type>AI_XOR2</type>
<position>-264,-68.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>505 </input>
<output>
<ID>OUT</ID>511 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>332</ID>
<type>AI_XOR2</type>
<position>-264,-72.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>504 </input>
<output>
<ID>OUT</ID>512 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>333</ID>
<type>AI_XOR2</type>
<position>-264,-76.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>503 </input>
<output>
<ID>OUT</ID>513 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>334</ID>
<type>AI_XOR2</type>
<position>-264,-80.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>514 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>335</ID>
<type>DD_KEYPAD_HEX</type>
<position>-277,-37</position>
<output>
<ID>OUT_0</ID>501 </output>
<output>
<ID>OUT_1</ID>500 </output>
<output>
<ID>OUT_2</ID>499 </output>
<output>
<ID>OUT_3</ID>498 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>336</ID>
<type>AI_XOR2</type>
<position>-194,-66.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>491 </input>
<output>
<ID>OUT</ID>495 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>337</ID>
<type>AA_TOGGLE</type>
<position>-266,-10.5</position>
<output>
<ID>OUT_0</ID>445 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>338</ID>
<type>AI_XOR2</type>
<position>-194,-70.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>490 </input>
<output>
<ID>OUT</ID>496 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>339</ID>
<type>DD_KEYPAD_HEX</type>
<position>-303.5,-54</position>
<output>
<ID>OUT_0</ID>456 </output>
<output>
<ID>OUT_1</ID>457 </output>
<output>
<ID>OUT_2</ID>463 </output>
<output>
<ID>OUT_3</ID>464 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>340</ID>
<type>AI_XOR2</type>
<position>-194,-74.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>490 </input>
<output>
<ID>OUT</ID>497 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>AI_XOR2</type>
<position>-194,-78.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>494 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>342</ID>
<type>DD_KEYPAD_HEX</type>
<position>-278.5,-78</position>
<output>
<ID>OUT_0</ID>505 </output>
<output>
<ID>OUT_1</ID>504 </output>
<output>
<ID>OUT_2</ID>503 </output>
<output>
<ID>OUT_3</ID>502 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>343</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-245,-42.5</position>
<input>
<ID>IN_0</ID>456 </input>
<input>
<ID>IN_1</ID>457 </input>
<input>
<ID>IN_2</ID>463 </input>
<input>
<ID>IN_3</ID>464 </input>
<input>
<ID>IN_B_0</ID>507 </input>
<input>
<ID>IN_B_1</ID>508 </input>
<input>
<ID>IN_B_2</ID>509 </input>
<input>
<ID>IN_B_3</ID>510 </input>
<output>
<ID>OUT_0</ID>446 </output>
<output>
<ID>OUT_1</ID>448 </output>
<output>
<ID>OUT_2</ID>447 </output>
<output>
<ID>OUT_3</ID>449 </output>
<input>
<ID>carry_in</ID>493 </input>
<output>
<ID>carry_out</ID>467 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>344</ID>
<type>DD_KEYPAD_HEX</type>
<position>-303,-91.5</position>
<output>
<ID>OUT_0</ID>455 </output>
<output>
<ID>OUT_1</ID>454 </output>
<output>
<ID>OUT_2</ID>453 </output>
<output>
<ID>OUT_3</ID>452 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>345</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-245,-82.5</position>
<input>
<ID>IN_0</ID>455 </input>
<input>
<ID>IN_1</ID>454 </input>
<input>
<ID>IN_2</ID>453 </input>
<input>
<ID>IN_3</ID>452 </input>
<input>
<ID>IN_B_0</ID>511 </input>
<input>
<ID>IN_B_1</ID>512 </input>
<input>
<ID>IN_B_2</ID>513 </input>
<input>
<ID>IN_B_3</ID>514 </input>
<output>
<ID>OUT_0</ID>458 </output>
<output>
<ID>OUT_1</ID>460 </output>
<output>
<ID>OUT_2</ID>459 </output>
<output>
<ID>OUT_3</ID>461 </output>
<input>
<ID>carry_in</ID>525 </input>
<output>
<ID>carry_out</ID>506 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>346</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-186,-29.5</position>
<input>
<ID>IN_0</ID>486 </input>
<input>
<ID>IN_1</ID>485 </input>
<input>
<ID>IN_2</ID>484 </input>
<input>
<ID>IN_3</ID>487 </input>
<input>
<ID>IN_B_0</ID>446 </input>
<input>
<ID>IN_B_1</ID>448 </input>
<input>
<ID>IN_B_2</ID>447 </input>
<input>
<ID>IN_B_3</ID>449 </input>
<output>
<ID>OUT_0</ID>471 </output>
<output>
<ID>OUT_1</ID>470 </output>
<output>
<ID>OUT_2</ID>469 </output>
<output>
<ID>OUT_3</ID>468 </output>
<input>
<ID>carry_in</ID>493 </input>
<output>
<ID>carry_out</ID>479 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>347</ID>
<type>AI_XOR2</type>
<position>-263,-27.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>348</ID>
<type>AI_XOR2</type>
<position>-263,-31.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>500 </input>
<output>
<ID>OUT</ID>508 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>349</ID>
<type>AA_LABEL</type>
<position>-299,-31.5</position>
<gparam>LABEL_TEXT /</gparam>
<gparam>TEXT_HEIGHT 12</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>-212,-46</position>
<output>
<ID>A_less_B</ID>472 </output>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_3</ID>450 </input>
<input>
<ID>IN_B_0</ID>446 </input>
<input>
<ID>IN_B_1</ID>448 </input>
<input>
<ID>IN_B_2</ID>447 </input>
<input>
<ID>IN_B_3</ID>449 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>351</ID>
<type>EE_VDD</type>
<position>-222,-51</position>
<output>
<ID>OUT_0</ID>450 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>352</ID>
<type>EE_VDD</type>
<position>-221.5,-48</position>
<output>
<ID>OUT_0</ID>451 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>353</ID>
<type>AA_LABEL</type>
<position>-276,-10</position>
<gparam>LABEL_TEXT is minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>354</ID>
<type>AA_TOGGLE</type>
<position>-268,-10.5</position>
<output>
<ID>OUT_0</ID>444 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_LABEL</type>
<position>-254.5,-9.5</position>
<gparam>LABEL_TEXT pressd minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>356</ID>
<type>AI_XOR2</type>
<position>-267,-15.5</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>444 </input>
<output>
<ID>OUT</ID>493 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>AI_XOR2</type>
<position>-263,-35.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>499 </input>
<output>
<ID>OUT</ID>509 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>358</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-186,-66.5</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>496 </input>
<input>
<ID>IN_2</ID>497 </input>
<input>
<ID>IN_3</ID>494 </input>
<input>
<ID>IN_B_0</ID>458 </input>
<input>
<ID>IN_B_1</ID>460 </input>
<input>
<ID>IN_B_2</ID>459 </input>
<input>
<ID>IN_B_3</ID>461 </input>
<output>
<ID>OUT_0</ID>473 </output>
<output>
<ID>OUT_1</ID>474 </output>
<output>
<ID>OUT_2</ID>475 </output>
<output>
<ID>OUT_3</ID>476 </output>
<input>
<ID>carry_in</ID>479 </input>
<output>
<ID>carry_out</ID>520 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>359</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>-210,-81.5</position>
<output>
<ID>A_less_B</ID>523 </output>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_3</ID>462 </input>
<input>
<ID>IN_B_0</ID>458 </input>
<input>
<ID>IN_B_1</ID>460 </input>
<input>
<ID>IN_B_2</ID>459 </input>
<input>
<ID>IN_B_3</ID>461 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>360</ID>
<type>AI_XOR2</type>
<position>-263,-39.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>498 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>EE_VDD</type>
<position>-215.5,-86.5</position>
<output>
<ID>OUT_0</ID>462 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>362</ID>
<type>GA_LED</type>
<position>-162.5,-78</position>
<input>
<ID>N_in2</ID>465 </input>
<input>
<ID>N_in3</ID>482 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>363</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-164,-30</position>
<input>
<ID>IN_0</ID>471 </input>
<input>
<ID>IN_1</ID>470 </input>
<input>
<ID>IN_2</ID>469 </input>
<input>
<ID>IN_3</ID>468 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>364</ID>
<type>AE_OR2</type>
<position>-206.5,-51</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>515 </input>
<output>
<ID>OUT</ID>483 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>365</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-162.5,-67</position>
<input>
<ID>IN_0</ID>473 </input>
<input>
<ID>IN_1</ID>474 </input>
<input>
<ID>IN_2</ID>475 </input>
<input>
<ID>IN_3</ID>476 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>366</ID>
<type>AE_OR2</type>
<position>-203.5,-97.5</position>
<input>
<ID>IN_0</ID>523 </input>
<input>
<ID>IN_1</ID>506 </input>
<output>
<ID>OUT</ID>518 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>367</ID>
<type>AI_XOR2</type>
<position>-217,-83.5</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>479 </input>
<output>
<ID>OUT</ID>517 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>368</ID>
<type>EE_VDD</type>
<position>-221,-82.5</position>
<output>
<ID>OUT_0</ID>480 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>369</ID>
<type>GA_LED</type>
<position>-162.5,-80</position>
<input>
<ID>N_in0</ID>524 </input>
<input>
<ID>N_in2</ID>466 </input>
<input>
<ID>N_in3</ID>465 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>370</ID>
<type>GA_LED</type>
<position>-162.5,-82</position>
<input>
<ID>N_in0</ID>478 </input>
<input>
<ID>N_in2</ID>478 </input>
<input>
<ID>N_in3</ID>466 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>371</ID>
<type>GA_LED</type>
<position>-162.5,-84</position>
<input>
<ID>N_in1</ID>524 </input>
<input>
<ID>N_in3</ID>478 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>372</ID>
<type>AA_AND2</type>
<position>-247,-13</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>445 </input>
<output>
<ID>OUT</ID>482 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>373</ID>
<type>AI_XOR2</type>
<position>-194.5,-30.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>488 </input>
<output>
<ID>OUT</ID>486 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>AI_XOR2</type>
<position>-194.5,-34.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>483 </input>
<output>
<ID>OUT</ID>485 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>AI_XOR2</type>
<position>-194.5,-38.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>483 </input>
<output>
<ID>OUT</ID>484 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>376</ID>
<type>AI_XOR2</type>
<position>-194.5,-42.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>489 </input>
<output>
<ID>OUT</ID>487 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>377</ID>
<type>AI_XOR2</type>
<position>-234,-56</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>467 </input>
<output>
<ID>OUT</ID>515 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>378</ID>
<type>AI_XOR2</type>
<position>-199.5,-92.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>518 </input>
<output>
<ID>OUT</ID>490 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>FF_GND</type>
<position>-198.5,-31.5</position>
<output>
<ID>OUT_0</ID>488 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>380</ID>
<type>FF_GND</type>
<position>-198.5,-43.5</position>
<output>
<ID>OUT_0</ID>489 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>381</ID>
<type>FF_GND</type>
<position>-198,-67.5</position>
<output>
<ID>OUT_0</ID>491 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>382</ID>
<type>AE_SMALL_INVERTER</type>
<position>510,1</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>383</ID>
<type>AE_SMALL_INVERTER</type>
<position>509.5,18</position>
<input>
<ID>IN_0</ID>261 </input>
<output>
<ID>OUT_0</ID>768 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>384</ID>
<type>AE_SMALL_INVERTER</type>
<position>510,35</position>
<input>
<ID>IN_0</ID>261 </input>
<output>
<ID>OUT_0</ID>769 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>385</ID>
<type>GA_LED</type>
<position>-172,-78.5</position>
<input>
<ID>N_in3</ID>520 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>386</ID>
<type>AE_OR2</type>
<position>-245,-70</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>467 </input>
<output>
<ID>OUT</ID>525 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>387</ID>
<type>AI_XOR2</type>
<position>326,-63</position>
<input>
<ID>IN_0</ID>530 </input>
<input>
<ID>IN_1</ID>545 </input>
<output>
<ID>OUT</ID>534 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>388</ID>
<type>AI_XOR2</type>
<position>330,-63</position>
<input>
<ID>IN_0</ID>530 </input>
<input>
<ID>IN_1</ID>544 </input>
<output>
<ID>OUT</ID>533 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>769</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,32.5,510,33</points>
<connection>
<GID>384</GID>
<name>OUT_0</name></connection>
<intersection>32.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>511,32,511,32.5</points>
<connection>
<GID>312</GID>
<name>shift_enable</name></connection>
<intersection>32.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>510,32.5,511,32.5</points>
<intersection>510 0</intersection>
<intersection>511 1</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-9,61,-8.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-8.5,79,-8.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-10.5,63,-9</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-10.5,79,-10.5</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-36,80,-36</points>
<connection>
<GID>14</GID>
<name>OUT_2</name></connection>
<connection>
<GID>22</GID>
<name>IN_B_2</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-35,80,-35</points>
<connection>
<GID>14</GID>
<name>OUT_1</name></connection>
<connection>
<GID>22</GID>
<name>IN_B_1</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-41.5,226.5,-39</points>
<intersection>-41.5 3</intersection>
<intersection>-39 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-41.5,226.5,-41.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-39,236,-39</points>
<connection>
<GID>66</GID>
<name>IN_B_0</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-40,226.5,-39.5</points>
<intersection>-40 6</intersection>
<intersection>-39.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>217,-39.5,226.5,-39.5</points>
<connection>
<GID>62</GID>
<name>OUT_1</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>226.5,-40,236,-40</points>
<connection>
<GID>66</GID>
<name>IN_B_1</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-41,226.5,-37.5</points>
<intersection>-41 4</intersection>
<intersection>-37.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-37.5,226.5,-37.5</points>
<connection>
<GID>62</GID>
<name>OUT_2</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-41,236,-41</points>
<connection>
<GID>66</GID>
<name>IN_B_2</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-42,226.5,-35.5</points>
<intersection>-42 4</intersection>
<intersection>-35.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-35.5,226.5,-35.5</points>
<connection>
<GID>62</GID>
<name>OUT_3</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-42,236,-42</points>
<connection>
<GID>66</GID>
<name>IN_B_3</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-42.5,273,-42.5</points>
<connection>
<GID>75</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>252.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>252.5,-42.5,252.5,-26</points>
<intersection>-42.5 1</intersection>
<intersection>-26 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>252.5,-26,285,-26</points>
<connection>
<GID>67</GID>
<name>IN_B_0</name></connection>
<intersection>252.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-44.5,273,-44.5</points>
<connection>
<GID>75</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>66</GID>
<name>OUT_2</name></connection>
<intersection>254.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>254.5,-44.5,254.5,-28</points>
<intersection>-44.5 1</intersection>
<intersection>-28 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>254.5,-28,285,-28</points>
<connection>
<GID>67</GID>
<name>IN_B_2</name></connection>
<intersection>254.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-43.5,273,-43.5</points>
<connection>
<GID>75</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>66</GID>
<name>OUT_1</name></connection>
<intersection>253.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>253.5,-43.5,253.5,-27</points>
<intersection>-43.5 1</intersection>
<intersection>-27 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>253.5,-27,285,-27</points>
<connection>
<GID>67</GID>
<name>IN_B_1</name></connection>
<intersection>253.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-45.5,273,-45.5</points>
<connection>
<GID>75</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>66</GID>
<name>OUT_3</name></connection>
<intersection>256 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>256,-45.5,256,-29</points>
<intersection>-45.5 1</intersection>
<intersection>-29 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>256,-29,285,-29</points>
<connection>
<GID>67</GID>
<name>IN_B_3</name></connection>
<intersection>256 6</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>268,-52.5,273,-52.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<connection>
<GID>75</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>268.5,-49.5,273,-49.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<connection>
<GID>75</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-49,213,-47.5</points>
<intersection>-49 4</intersection>
<intersection>-47.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>190.5,-47.5,213,-47.5</points>
<connection>
<GID>64</GID>
<name>OUT_3</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>213,-49,236,-49</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-49.5,213,-48</points>
<intersection>-49.5 3</intersection>
<intersection>-48 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>190.5,-49.5,213,-49.5</points>
<connection>
<GID>64</GID>
<name>OUT_2</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>213,-48,236,-48</points>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-51.5,213,-47</points>
<intersection>-51.5 3</intersection>
<intersection>-47 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>190.5,-51.5,213,-51.5</points>
<connection>
<GID>64</GID>
<name>OUT_1</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>213,-47,236,-47</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-53.5,213,-46</points>
<intersection>-53.5 3</intersection>
<intersection>-46 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>190.5,-53.5,213,-53.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>213,-46,236,-46</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>283.5,-50,283.5,-34</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>-35 30</intersection>
<intersection>-34 31</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>283.5,-35,285,-35</points>
<connection>
<GID>67</GID>
<name>IN_2</name></connection>
<intersection>283.5 2</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>283.5,-34,285,-34</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>283.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-78,226.5,-74.5</points>
<intersection>-78 3</intersection>
<intersection>-74.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217.5,-78,226.5,-78</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-74.5,236,-74.5</points>
<connection>
<GID>85</GID>
<name>IN_B_0</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-76,226.5,-75.5</points>
<intersection>-76 7</intersection>
<intersection>-75.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>217.5,-76,226.5,-76</points>
<connection>
<GID>83</GID>
<name>OUT_1</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>226.5,-75.5,236,-75.5</points>
<connection>
<GID>85</GID>
<name>IN_B_1</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-76.5,226.5,-74</points>
<intersection>-76.5 4</intersection>
<intersection>-74 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217.5,-74,226.5,-74</points>
<connection>
<GID>83</GID>
<name>OUT_2</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-76.5,236,-76.5</points>
<connection>
<GID>85</GID>
<name>IN_B_2</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-77.5,226.5,-72</points>
<intersection>-77.5 4</intersection>
<intersection>-72 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217.5,-72,226.5,-72</points>
<connection>
<GID>83</GID>
<name>OUT_3</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-77.5,236,-77.5</points>
<connection>
<GID>85</GID>
<name>IN_B_3</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-37.5,113,-37.5</points>
<connection>
<GID>37</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>92.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>92.5,-37.5,92.5,-21</points>
<intersection>-37.5 1</intersection>
<intersection>-21 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>92.5,-21,139,-21</points>
<connection>
<GID>27</GID>
<name>IN_B_0</name></connection>
<intersection>92.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-39.5,113,-39.5</points>
<connection>
<GID>37</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>22</GID>
<name>OUT_2</name></connection>
<intersection>94.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>94.5,-39.5,94.5,-23</points>
<intersection>-39.5 1</intersection>
<intersection>-23 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>94.5,-23,139,-23</points>
<connection>
<GID>27</GID>
<name>IN_B_2</name></connection>
<intersection>94.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-38.5,113,-38.5</points>
<connection>
<GID>37</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>22</GID>
<name>OUT_1</name></connection>
<intersection>93.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>93.5,-38.5,93.5,-22</points>
<intersection>-38.5 1</intersection>
<intersection>-22 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>93.5,-22,139,-22</points>
<connection>
<GID>27</GID>
<name>IN_B_1</name></connection>
<intersection>93.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-40.5,113,-40.5</points>
<connection>
<GID>37</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>22</GID>
<name>OUT_3</name></connection>
<intersection>96 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>96,-40.5,96,-24</points>
<intersection>-40.5 1</intersection>
<intersection>-24 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>96,-24,139,-24</points>
<connection>
<GID>27</GID>
<name>IN_B_3</name></connection>
<intersection>96 6</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-47.5,113,-47.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108.5,-44.5,113,-44.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-78,276.5,-78</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<connection>
<GID>92</GID>
<name>IN_B_0</name></connection>
<intersection>255 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>255,-78,255,-63</points>
<intersection>-78 1</intersection>
<intersection>-63 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>255,-63,287.5,-63</points>
<connection>
<GID>86</GID>
<name>IN_B_0</name></connection>
<intersection>255 6</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-37,80,-37</points>
<connection>
<GID>14</GID>
<name>OUT_3</name></connection>
<connection>
<GID>22</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-34,80,-34</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<connection>
<GID>22</GID>
<name>IN_B_0</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-92.5,80,-92.5</points>
<intersection>31 5</intersection>
<intersection>80 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>31,-92.5,31,-85</points>
<connection>
<GID>216</GID>
<name>OUT_3</name></connection>
<intersection>-92.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>80,-92.5,80,-84</points>
<connection>
<GID>217</GID>
<name>IN_3</name></connection>
<intersection>-92.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-92.5,80,-83</points>
<connection>
<GID>217</GID>
<name>IN_2</name></connection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-92.5,80,-92.5</points>
<intersection>31 3</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-92.5,31,-87</points>
<connection>
<GID>216</GID>
<name>OUT_2</name></connection>
<intersection>-92.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-36,69.5,-33.5</points>
<intersection>-36 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-33.5,72,-33.5</points>
<connection>
<GID>14</GID>
<name>IN_B_3</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-36,69.5,-36</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-80,276.5,-80</points>
<connection>
<GID>85</GID>
<name>OUT_2</name></connection>
<connection>
<GID>92</GID>
<name>IN_B_2</name></connection>
<intersection>257 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>257,-80,257,-65</points>
<intersection>-80 1</intersection>
<intersection>-65 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>257,-65,287.5,-65</points>
<connection>
<GID>86</GID>
<name>IN_B_2</name></connection>
<intersection>257 6</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-79,276.5,-79</points>
<connection>
<GID>85</GID>
<name>OUT_1</name></connection>
<connection>
<GID>92</GID>
<name>IN_B_1</name></connection>
<intersection>256 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>256,-79,256,-64</points>
<intersection>-79 1</intersection>
<intersection>-64 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>256,-64,287.5,-64</points>
<connection>
<GID>86</GID>
<name>IN_B_1</name></connection>
<intersection>256 8</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-81,276.5,-81</points>
<connection>
<GID>85</GID>
<name>OUT_3</name></connection>
<connection>
<GID>92</GID>
<name>IN_B_3</name></connection>
<intersection>258.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>258.5,-81,258.5,-66</points>
<intersection>-81 1</intersection>
<intersection>-66 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>258.5,-66,287.5,-66</points>
<connection>
<GID>86</GID>
<name>IN_B_3</name></connection>
<intersection>258.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>276.5,-88,276.5,-88</points>
<connection>
<GID>92</GID>
<name>IN_3</name></connection>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-92.5,80,-82</points>
<connection>
<GID>217</GID>
<name>IN_1</name></connection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-92.5,80,-92.5</points>
<intersection>31 3</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-92.5,31,-89</points>
<connection>
<GID>216</GID>
<name>OUT_1</name></connection>
<intersection>-92.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-92.5,80,-81</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-92.5,80,-92.5</points>
<intersection>31 3</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-92.5,31,-91</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>-92.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-53,80,-41</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-53,80,-53</points>
<intersection>30.5 3</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-53,30.5,-50</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>-53 2</intersection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-51.5,80,-42</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-51.5,80,-51.5</points>
<intersection>30.5 3</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-51.5,30.5,-48</points>
<connection>
<GID>19</GID>
<name>OUT_1</name></connection>
<intersection>-51.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88.5,-73,116.5,-73</points>
<connection>
<GID>55</GID>
<name>IN_B_0</name></connection>
<intersection>88.5 9</intersection>
<intersection>95 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>95,-73,95,-58</points>
<intersection>-73 1</intersection>
<intersection>-58 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>95,-58,139,-58</points>
<connection>
<GID>54</GID>
<name>IN_B_0</name></connection>
<intersection>95 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>88.5,-77.5,88.5,-73</points>
<intersection>-77.5 12</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>88,-77.5,88.5,-77.5</points>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<intersection>88.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91,-75,116.5,-75</points>
<connection>
<GID>55</GID>
<name>IN_B_2</name></connection>
<intersection>91 8</intersection>
<intersection>97 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>97,-75,97,-60</points>
<intersection>-75 1</intersection>
<intersection>-60 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>97,-60,139,-60</points>
<connection>
<GID>54</GID>
<name>IN_B_2</name></connection>
<intersection>97 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>91,-79.5,91,-75</points>
<intersection>-79.5 9</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>88,-79.5,91,-79.5</points>
<connection>
<GID>217</GID>
<name>OUT_2</name></connection>
<intersection>91 8</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,-74,116.5,-74</points>
<connection>
<GID>55</GID>
<name>IN_B_1</name></connection>
<intersection>90 10</intersection>
<intersection>96 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>96,-74,96,-59</points>
<intersection>-74 1</intersection>
<intersection>-59 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>96,-59,139,-59</points>
<connection>
<GID>54</GID>
<name>IN_B_1</name></connection>
<intersection>96 8</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>90,-78.5,90,-74</points>
<intersection>-78.5 14</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>88,-78.5,90,-78.5</points>
<connection>
<GID>217</GID>
<name>OUT_1</name></connection>
<intersection>90 10</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-76,116.5,-76</points>
<connection>
<GID>55</GID>
<name>IN_B_3</name></connection>
<intersection>93.5 8</intersection>
<intersection>98.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>98.5,-76,98.5,-61</points>
<intersection>-76 1</intersection>
<intersection>-61 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>98.5,-61,139,-61</points>
<connection>
<GID>54</GID>
<name>IN_B_3</name></connection>
<intersection>98.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>93.5,-80.5,93.5,-76</points>
<intersection>-80.5 9</intersection>
<intersection>-76 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>88,-80.5,93.5,-80.5</points>
<connection>
<GID>217</GID>
<name>OUT_3</name></connection>
<intersection>93.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>116.5,-83,116.5,-83</points>
<connection>
<GID>55</GID>
<name>IN_3</name></connection>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-50.5,79.5,-43</points>
<intersection>-50.5 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-50.5,79.5,-50.5</points>
<intersection>30.5 3</intersection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79.5,-43,80,-43</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>79.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-50.5,30.5,-46</points>
<connection>
<GID>19</GID>
<name>OUT_2</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-49.5,80,-49.5</points>
<intersection>30.5 3</intersection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-49.5,80,-44</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-49.5,30.5,-44</points>
<connection>
<GID>19</GID>
<name>OUT_3</name></connection>
<intersection>-49.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>166.5,-75.5,166.5,-75.5</points>
<connection>
<GID>63</GID>
<name>N_in2</name></connection>
<connection>
<GID>81</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>166.5,-77.5,166.5,-77.5</points>
<connection>
<GID>81</GID>
<name>N_in2</name></connection>
<connection>
<GID>129</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-32.5,72,-32.5</points>
<connection>
<GID>14</GID>
<name>IN_B_2</name></connection>
<intersection>69 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>69,-32.5,69,-32</points>
<connection>
<GID>199</GID>
<name>OUT</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-84.5,214.5,-84</points>
<intersection>-84.5 5</intersection>
<intersection>-84 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>193,-84,214.5,-84</points>
<connection>
<GID>84</GID>
<name>OUT_3</name></connection>
<intersection>214.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>214.5,-84.5,236,-84.5</points>
<connection>
<GID>85</GID>
<name>IN_3</name></connection>
<intersection>214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-86,214.5,-83.5</points>
<intersection>-86 3</intersection>
<intersection>-83.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>193,-86,214.5,-86</points>
<connection>
<GID>84</GID>
<name>OUT_2</name></connection>
<intersection>214.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>214.5,-83.5,236,-83.5</points>
<connection>
<GID>85</GID>
<name>IN_2</name></connection>
<intersection>214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-88,214.5,-82.5</points>
<intersection>-88 3</intersection>
<intersection>-82.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>193,-88,214.5,-88</points>
<connection>
<GID>84</GID>
<name>OUT_1</name></connection>
<intersection>214.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>214.5,-82.5,236,-82.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-71,83,-47</points>
<connection>
<GID>22</GID>
<name>carry_out</name></connection>
<connection>
<GID>217</GID>
<name>carry_in</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-53.5,123.5,-53.5</points>
<intersection>83 0</intersection>
<intersection>123.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123.5,-53.5,123.5,-50.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>-53.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-90,214.5,-81.5</points>
<intersection>-90 3</intersection>
<intersection>-81.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>193,-90,214.5,-90</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>214.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>214.5,-81.5,236,-81.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-27.5,162,-24.5</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-27.5,162,-27.5</points>
<connection>
<GID>27</GID>
<name>OUT_3</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-26.5,162,-25.5</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-26.5,162,-26.5</points>
<connection>
<GID>27</GID>
<name>OUT_2</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>162,-26.5,162,-25.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>-25.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>147,-25.5,162,-25.5</points>
<connection>
<GID>27</GID>
<name>OUT_1</name></connection>
<intersection>162 3</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-27.5,162,-24.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-24.5,162,-24.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>289,-94.5,289,-77.5</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>-77.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>286.5,-77.5,289,-77.5</points>
<intersection>286.5 10</intersection>
<intersection>289 2</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>286.5,-77.5,286.5,-71</points>
<intersection>-77.5 8</intersection>
<intersection>-72 12</intersection>
<intersection>-71 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>286.5,-71,287.5,-71</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>286.5 10</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>286.5,-72,287.5,-72</points>
<connection>
<GID>86</GID>
<name>IN_2</name></connection>
<intersection>286.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>119,-51,121.5,-51</points>
<intersection>119 6</intersection>
<intersection>121.5 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>119,-51,119,-50.5</points>
<connection>
<GID>37</GID>
<name>A_less_B</name></connection>
<intersection>-51 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>121.5,-51,121.5,-50.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>-51 2</intersection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-71.5,239,-52</points>
<connection>
<GID>66</GID>
<name>carry_out</name></connection>
<connection>
<GID>85</GID>
<name>carry_in</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,-58,284.5,-58</points>
<intersection>239 0</intersection>
<intersection>284.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>284.5,-58,284.5,-56</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>-58 1</intersection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295,-32.5,295,-29</points>
<intersection>-32.5 1</intersection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293,-32.5,295,-32.5</points>
<connection>
<GID>67</GID>
<name>OUT_3</name></connection>
<intersection>295 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295,-29,299,-29</points>
<connection>
<GID>114</GID>
<name>IN_3</name></connection>
<intersection>295 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-64.5,163.5,-61.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-61.5,163.5,-61.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-63.5,146.5,-62.5</points>
<intersection>-63.5 1</intersection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>146.5,-63.5,163.5,-63.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>146.5,-62.5,147,-62.5</points>
<connection>
<GID>54</GID>
<name>OUT_1</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-63.5,163.5,-62.5</points>
<connection>
<GID>73</GID>
<name>IN_2</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-63.5,163.5,-63.5</points>
<connection>
<GID>54</GID>
<name>OUT_2</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164,-64.5,164,-61.5</points>
<intersection>-64.5 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-64.5,164,-64.5</points>
<connection>
<GID>54</GID>
<name>OUT_3</name></connection>
<intersection>164 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163.5,-61.5,164,-61.5</points>
<connection>
<GID>73</GID>
<name>IN_3</name></connection>
<intersection>164 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-88.5,122.5,-86</points>
<connection>
<GID>55</GID>
<name>A_less_B</name></connection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-88.5,123,-88.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166,-79.5,166.5,-79.5</points>
<connection>
<GID>174</GID>
<name>N_in3</name></connection>
<connection>
<GID>129</GID>
<name>N_in2</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-79.5,166,-78.5</points>
<intersection>-79.5 1</intersection>
<intersection>-78.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>165.5,-78.5,166,-78.5</points>
<connection>
<GID>129</GID>
<name>N_in0</name></connection>
<intersection>166 4</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-55,142,-34</points>
<connection>
<GID>54</GID>
<name>carry_in</name></connection>
<connection>
<GID>27</GID>
<name>carry_out</name></connection>
<intersection>-54.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>104,-54.5,142,-54.5</points>
<intersection>104 9</intersection>
<intersection>142 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>104,-81,104,-54.5</points>
<intersection>-81 10</intersection>
<intersection>-54.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>104,-81,109,-81</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>104 9</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295,-31.5,295,-30</points>
<intersection>-31.5 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293,-31.5,295,-31.5</points>
<connection>
<GID>67</GID>
<name>OUT_2</name></connection>
<intersection>295 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295,-30,299,-30</points>
<connection>
<GID>114</GID>
<name>IN_2</name></connection>
<intersection>295 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-79,109,-79</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>293,-31,299,-31</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>293 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>293,-31,293,-30.5</points>
<connection>
<GID>67</GID>
<name>OUT_1</name></connection>
<intersection>-31 1</intersection></vsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296,-32,296,-29.5</points>
<intersection>-32 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293,-29.5,296,-29.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>296 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>296,-32,299,-32</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>296 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>279,-56,282.5,-56</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>279 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>279,-56,279,-55.5</points>
<connection>
<GID>75</GID>
<name>A_less_B</name></connection>
<intersection>-56 2</intersection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>115,-80,116.5,-80</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>78</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-69.5,298,-66.5</points>
<intersection>-69.5 2</intersection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-66.5,298,-66.5</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>298 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>298,-69.5,300.5,-69.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>298 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-68.5,298,-67.5</points>
<intersection>-68.5 1</intersection>
<intersection>-67.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>298,-68.5,300.5,-68.5</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>298 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295.5,-67.5,298,-67.5</points>
<connection>
<GID>86</GID>
<name>OUT_1</name></connection>
<intersection>298 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-68.5,298,-67.5</points>
<intersection>-68.5 1</intersection>
<intersection>-67.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-68.5,298,-68.5</points>
<connection>
<GID>86</GID>
<name>OUT_2</name></connection>
<intersection>298 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>298,-67.5,300.5,-67.5</points>
<connection>
<GID>120</GID>
<name>IN_2</name></connection>
<intersection>298 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-69.5,298,-66.5</points>
<intersection>-69.5 1</intersection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-69.5,298,-69.5</points>
<connection>
<GID>86</GID>
<name>OUT_3</name></connection>
<intersection>298 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>298,-66.5,300.5,-66.5</points>
<connection>
<GID>120</GID>
<name>IN_3</name></connection>
<intersection>298 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282.5,-93.5,282.5,-91</points>
<connection>
<GID>92</GID>
<name>A_less_B</name></connection>
<intersection>-93.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282.5,-93.5,283,-93.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>282.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-95.5,239,-87.5</points>
<connection>
<GID>85</GID>
<name>carry_out</name></connection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,-95.5,283,-95.5</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-60,288,-39</points>
<connection>
<GID>67</GID>
<name>carry_out</name></connection>
<intersection>-60 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>264,-60,290.5,-60</points>
<connection>
<GID>86</GID>
<name>carry_in</name></connection>
<intersection>264 6</intersection>
<intersection>288 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>264,-86,264,-60</points>
<intersection>-86 7</intersection>
<intersection>-60 3</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>264,-86,269,-86</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>264 6</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>269,-84,269,-84</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>275,-85,276.5,-85</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-73.5,172,-9.5</points>
<intersection>-73.5 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-9.5,172,-9.5</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>172 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,-73.5,172,-73.5</points>
<connection>
<GID>63</GID>
<name>N_in3</name></connection>
<intersection>172 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-44.5,122.5,-32</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>-36 21</intersection>
<intersection>-32 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>122.5,-32,131.5,-32</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>122.5,-36,131.5,-36</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-35,138.5,-30</points>
<intersection>-35 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-30,139,-30</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-35,138.5,-35</points>
<connection>
<GID>191</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-31,138,-29</points>
<intersection>-31 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-29,139,-29</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-31,138,-31</points>
<connection>
<GID>190</GID>
<name>OUT</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-28,138,-27</points>
<intersection>-28 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-28,139,-28</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-27,138,-27</points>
<connection>
<GID>189</GID>
<name>OUT</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-39,139,-31</points>
<connection>
<GID>27</GID>
<name>IN_3</name></connection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-39,139,-39</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-31.5,69.5,-28</points>
<intersection>-31.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-31.5,72,-31.5</points>
<connection>
<GID>14</GID>
<name>IN_B_1</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-28,69.5,-28</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-28,131.5,-28</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-40,131.5,-40</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-89.5,129,-68</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>-72 21</intersection>
<intersection>-68 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>129,-68,132,-68</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>129,-72,132,-72</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-64,132,-64</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<connection>
<GID>210</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-76,132,-76</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<connection>
<GID>213</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-30.5,69.5,-24</points>
<intersection>-30.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-24,69.5,-24</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-30.5,72,-30.5</points>
<connection>
<GID>14</GID>
<name>IN_B_0</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-80.5,62,-15</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>-80.5 136</intersection>
<intersection>-40.5 31</intersection>
<intersection>-35 101</intersection>
<intersection>-31 39</intersection>
<intersection>-27 29</intersection>
<intersection>-23 28</intersection>
<intersection>-15 30</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>62,-23,63,-23</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>62,-27,63,-27</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>62,-15,142,-15</points>
<intersection>62 0</intersection>
<intersection>127.5 37</intersection>
<intersection>142 226</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>62,-40.5,75,-40.5</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<intersection>62 0</intersection>
<intersection>70.5 224</intersection>
<intersection>75 222</intersection></hsegment>
<vsegment>
<ID>37</ID>
<points>127.5,-74,127.5,-15</points>
<intersection>-74 90</intersection>
<intersection>-70 98</intersection>
<intersection>-66 95</intersection>
<intersection>-62 96</intersection>
<intersection>-38 40</intersection>
<intersection>-34 48</intersection>
<intersection>-30 45</intersection>
<intersection>-26 228</intersection>
<intersection>-15 30</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>62,-31,63,-31</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>127.5,-38,131.5,-38</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>127.5,-30,131.5,-30</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>127.5,-34,131.5,-34</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>90</ID>
<points>127.5,-74,132,-74</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>95</ID>
<points>127.5,-66,132,-66</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>96</ID>
<points>127.5,-62,132,-62</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>98</ID>
<points>127.5,-70,132,-70</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>101</ID>
<points>62,-35,63,-35</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>136</ID>
<points>62,-80.5,72,-80.5</points>
<connection>
<GID>41</GID>
<name>IN_3</name></connection>
<intersection>62 0</intersection>
<intersection>71.5 218</intersection></hsegment>
<vsegment>
<ID>218</ID>
<points>71.5,-80.5,71.5,-77.5</points>
<intersection>-80.5 136</intersection>
<intersection>-77.5 221</intersection></vsegment>
<hsegment>
<ID>221</ID>
<points>71.5,-77.5,75,-77.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>71.5 218</intersection>
<intersection>75 223</intersection></hsegment>
<vsegment>
<ID>222</ID>
<points>75,-40.5,75,-27.5</points>
<connection>
<GID>14</GID>
<name>carry_in</name></connection>
<intersection>-40.5 31</intersection></vsegment>
<vsegment>
<ID>223</ID>
<points>75,-77.5,75,-67.5</points>
<connection>
<GID>41</GID>
<name>carry_in</name></connection>
<intersection>-77.5 221</intersection></vsegment>
<vsegment>
<ID>224</ID>
<points>70.5,-40.5,70.5,-37.5</points>
<intersection>-40.5 31</intersection>
<intersection>-37.5 225</intersection></vsegment>
<hsegment>
<ID>225</ID>
<points>70.5,-37.5,72,-37.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>70.5 224</intersection></hsegment>
<vsegment>
<ID>226</ID>
<points>142,-18,142,-15</points>
<connection>
<GID>27</GID>
<name>carry_in</name></connection>
<intersection>-15 30</intersection></vsegment>
<hsegment>
<ID>228</ID>
<points>127.5,-26,131.5,-26</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>518,-18,518,33</points>
<connection>
<GID>672</GID>
<name>OUT_0</name></connection>
<intersection>3 9</intersection>
<intersection>16.5 4</intersection>
<intersection>33 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>511,16.5,518,16.5</points>
<intersection>511 7</intersection>
<intersection>518 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>512,33,518,33</points>
<intersection>512 8</intersection>
<intersection>517.5 13</intersection>
<intersection>518 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>511,15,511,19</points>
<connection>
<GID>313</GID>
<name>load</name></connection>
<intersection>16.5 4</intersection>
<intersection>19 16</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>512,32,512,33</points>
<connection>
<GID>312</GID>
<name>load</name></connection>
<intersection>33 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>510,3,518,3</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>511 11</intersection>
<intersection>518 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>511,-1,511,3</points>
<connection>
<GID>325</GID>
<name>load</name></connection>
<intersection>3 9</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>517.5,33,517.5,37.5</points>
<intersection>33 6</intersection>
<intersection>37.5 20</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>509.5,19,511,19</points>
<intersection>509.5 21</intersection>
<intersection>511 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>510,37.5,517.5,37.5</points>
<intersection>510 22</intersection>
<intersection>517.5 13</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>509.5,19,509.5,20</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>19 16</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>510,37,510,37.5</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>37.5 20</intersection></vsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-76,80,-76</points>
<connection>
<GID>41</GID>
<name>OUT_2</name></connection>
<connection>
<GID>217</GID>
<name>IN_B_2</name></connection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-74,80,-74</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<connection>
<GID>217</GID>
<name>IN_B_0</name></connection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-75,80,-75</points>
<connection>
<GID>41</GID>
<name>OUT_1</name></connection>
<connection>
<GID>217</GID>
<name>IN_B_1</name></connection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-75,139,-68</points>
<connection>
<GID>54</GID>
<name>IN_3</name></connection>
<intersection>-75 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138,-75,139,-75</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-77,80,-77</points>
<connection>
<GID>41</GID>
<name>OUT_3</name></connection>
<connection>
<GID>217</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-65,138.5,-63</points>
<intersection>-65 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-65,139,-65</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-63,138.5,-63</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-67,138,-66</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-66,139,-66</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-71,138.5,-67</points>
<intersection>-71 4</intersection>
<intersection>-67 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>138.5,-67,139,-67</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>138,-71,138.5,-71</points>
<connection>
<GID>212</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-37,61,-30.5</points>
<intersection>-37 5</intersection>
<intersection>-30.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>57,-30.5,61,-30.5</points>
<connection>
<GID>17</GID>
<name>OUT_3</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61,-37,63,-37</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-33,61,-32.5</points>
<intersection>-33 5</intersection>
<intersection>-32.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>57,-32.5,61,-32.5</points>
<connection>
<GID>17</GID>
<name>OUT_2</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61,-33,63,-33</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-34.5,61,-29</points>
<intersection>-34.5 4</intersection>
<intersection>-29 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>57,-34.5,61,-34.5</points>
<connection>
<GID>17</GID>
<name>OUT_1</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61,-29,63,-29</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-36.5,61,-25</points>
<intersection>-36.5 4</intersection>
<intersection>-25 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>57,-36.5,61,-36.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61,-25,63,-25</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-70.5,70,-65</points>
<intersection>-70.5 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-70.5,72,-70.5</points>
<connection>
<GID>41</GID>
<name>IN_B_0</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-65,70,-65</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393.5,-11.5,393.5,-4</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<intersection>-11.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>384.5,-11.5,393.5,-11.5</points>
<connection>
<GID>228</GID>
<name>IN_B_0</name></connection>
<intersection>393.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>383.5,-11.5,383.5,-7.5</points>
<connection>
<GID>228</GID>
<name>IN_B_1</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>389.5,-7.5,389.5,-4</points>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>383.5,-7.5,389.5,-7.5</points>
<intersection>383.5 0</intersection>
<intersection>389.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>382.5,-11.5,382.5,-4</points>
<connection>
<GID>228</GID>
<name>IN_B_2</name></connection>
<intersection>-4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>382.5,-4,385.5,-4</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<intersection>382.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-71.5,69.5,-69</points>
<intersection>-71.5 2</intersection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-69,69.5,-69</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-71.5,72,-71.5</points>
<connection>
<GID>41</GID>
<name>IN_B_1</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381.5,-11.5,381.5,-4</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<connection>
<GID>228</GID>
<name>IN_B_3</name></connection></vsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-73,70,-72.5</points>
<intersection>-73 1</intersection>
<intersection>-72.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-73,70,-73</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-72.5,72,-72.5</points>
<connection>
<GID>41</GID>
<name>IN_B_2</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-77,70,-73.5</points>
<intersection>-77 1</intersection>
<intersection>-73.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-77,70,-77</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-73.5,72,-73.5</points>
<connection>
<GID>41</GID>
<name>IN_B_3</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-10.5,-106.5,-10</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-106.5,-10,-88.5,-10</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-104.5,-12,-104.5,-10.5</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-104.5,-12,-88.5,-12</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>-104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79.5,-39,-54.5,-39</points>
<connection>
<GID>252</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<intersection>-75 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-75,-39,-75,-22.5</points>
<intersection>-39 1</intersection>
<intersection>-22.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-75,-22.5,-28.5,-22.5</points>
<connection>
<GID>242</GID>
<name>IN_B_0</name></connection>
<intersection>-75 6</intersection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-78,60,-71.5</points>
<intersection>-78 3</intersection>
<intersection>-71.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>60,-78,62,-78</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>55.5,-71.5,60,-71.5</points>
<connection>
<GID>214</GID>
<name>OUT_3</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-74,60,-73.5</points>
<intersection>-74 3</intersection>
<intersection>-73.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>60,-74,62,-74</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>55.5,-73.5,60,-73.5</points>
<connection>
<GID>214</GID>
<name>OUT_2</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-75.5,60,-70</points>
<intersection>-75.5 4</intersection>
<intersection>-70 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>60,-70,62,-70</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>55.5,-75.5,60,-75.5</points>
<connection>
<GID>214</GID>
<name>OUT_1</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-77.5,60,-66</points>
<intersection>-77.5 4</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>60,-66,62,-66</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>55.5,-77.5,60,-77.5</points>
<connection>
<GID>214</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>343,4.5,402.5,4.5</points>
<intersection>343 18</intersection>
<intersection>345 21</intersection>
<intersection>351 25</intersection>
<intersection>355 24</intersection>
<intersection>359 23</intersection>
<intersection>363 22</intersection>
<intersection>374.5 5</intersection>
<intersection>376.5 8</intersection>
<intersection>382.5 26</intersection>
<intersection>386.5 27</intersection>
<intersection>390.5 28</intersection>
<intersection>394.5 29</intersection>
<intersection>402.5 9</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>374.5,-11.5,374.5,4.5</points>
<connection>
<GID>228</GID>
<name>IN_3</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>376.5,-11.5,376.5,4.5</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>402.5,4.5,402.5,36.5</points>
<intersection>4.5 1</intersection>
<intersection>36.5 11</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>365.5,36.5,365.5,37.5</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>36.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>363,36.5,402.5,36.5</points>
<connection>
<GID>259</GID>
<name>nQ</name></connection>
<intersection>365.5 10</intersection>
<intersection>402.5 9</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>343,-11.5,343,4.5</points>
<connection>
<GID>282</GID>
<name>IN_3</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>345,-11.5,345,4.5</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>363,2,363,4.5</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>359,2,359,4.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>355,2,355,4.5</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>351,2,351,4.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>382.5,2,382.5,4.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>386.5,2,386.5,4.5</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>390.5,2,390.5,4.5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>394.5,2,394.5,4.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79.5,-41,-54.5,-41</points>
<connection>
<GID>252</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>236</GID>
<name>OUT_2</name></connection>
<intersection>-73 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-73,-41,-73,-24.5</points>
<intersection>-41 1</intersection>
<intersection>-24.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-73,-24.5,-28.5,-24.5</points>
<connection>
<GID>242</GID>
<name>IN_B_2</name></connection>
<intersection>-73 6</intersection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79.5,-40,-54.5,-40</points>
<connection>
<GID>252</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>236</GID>
<name>OUT_1</name></connection>
<intersection>-74 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-74,-40,-74,-23.5</points>
<intersection>-40 1</intersection>
<intersection>-23.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-74,-23.5,-28.5,-23.5</points>
<connection>
<GID>242</GID>
<name>IN_B_1</name></connection>
<intersection>-74 8</intersection></hsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379,-22,379,-19.5</points>
<connection>
<GID>228</GID>
<name>OUT_2</name></connection>
<intersection>-22 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>373.5,-22,379,-22</points>
<intersection>373.5 16</intersection>
<intersection>379 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>373.5,-25,373.5,-22</points>
<connection>
<GID>241</GID>
<name>IN_B_2</name></connection>
<intersection>-22 5</intersection></vsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-90.5,83,-87</points>
<connection>
<GID>217</GID>
<name>carry_out</name></connection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-90.5,123,-90.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381,-25,381,-19.5</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>-25 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>375.5,-25,381,-25</points>
<connection>
<GID>241</GID>
<name>IN_B_0</name></connection>
<intersection>381 0</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372.5,-25,372.5,-19.5</points>
<connection>
<GID>241</GID>
<name>IN_B_3</name></connection>
<intersection>-19.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>372.5,-19.5,378,-19.5</points>
<connection>
<GID>228</GID>
<name>OUT_3</name></connection>
<intersection>372.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,-23,380,-19.5</points>
<connection>
<GID>228</GID>
<name>OUT_1</name></connection>
<intersection>-23 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>374.5,-23,380,-23</points>
<intersection>374.5 16</intersection>
<intersection>380 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>374.5,-25,374.5,-23</points>
<connection>
<GID>241</GID>
<name>IN_B_1</name></connection>
<intersection>-23 5</intersection></vsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79.5,-42,-54.5,-42</points>
<connection>
<GID>252</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>236</GID>
<name>OUT_3</name></connection>
<intersection>-71.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-71.5,-42,-71.5,-25.5</points>
<intersection>-42 1</intersection>
<intersection>-25.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-71.5,-25.5,-28.5,-25.5</points>
<connection>
<GID>242</GID>
<name>IN_B_3</name></connection>
<intersection>-71.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-49,-54.5,-49</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<connection>
<GID>252</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59,-46,-54.5,-46</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<connection>
<GID>252</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>523.5,-27,523.5,22</points>
<intersection>-27 16</intersection>
<intersection>-23 4</intersection>
<intersection>5 3</intersection>
<intersection>22 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>511,5,523.5,5</points>
<connection>
<GID>313</GID>
<name>clock</name></connection>
<intersection>523.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>495.5,-23,523.5,-23</points>
<connection>
<GID>670</GID>
<name>CLK</name></connection>
<intersection>511 7</intersection>
<intersection>523.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>512,22,523.5,22</points>
<connection>
<GID>312</GID>
<name>clock</name></connection>
<intersection>523.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>511,-23,511,-11</points>
<connection>
<GID>325</GID>
<name>clock</name></connection>
<intersection>-23 4</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>523.5,-27,533,-27</points>
<connection>
<GID>311</GID>
<name>clock</name></connection>
<intersection>523.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>508.5,-1,508.5,5</points>
<connection>
<GID>325</GID>
<name>carry_in</name></connection>
<connection>
<GID>313</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,21.5,366.5,40.5</points>
<connection>
<GID>264</GID>
<name>N_in2</name></connection>
<intersection>26.5 12</intersection>
<intersection>37.5 13</intersection>
<intersection>40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>363,40.5,366.5,40.5</points>
<connection>
<GID>259</GID>
<name>Q</name></connection>
<intersection>366.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>366.5,26.5,367.5,26.5</points>
<connection>
<GID>266</GID>
<name>N_in1</name></connection>
<intersection>366.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>366.5,37.5,367.5,37.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>366.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>357,36.5,357,40.5</points>
<connection>
<GID>259</GID>
<name>clock</name></connection>
<connection>
<GID>259</GID>
<name>K</name></connection>
<connection>
<GID>259</GID>
<name>J</name></connection>
<connection>
<GID>257</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,24.5,366.5,31.5</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>365.5,24.5,369.5,24.5</points>
<connection>
<GID>268</GID>
<name>N_in1</name></connection>
<connection>
<GID>261</GID>
<name>N_in1</name></connection>
<connection>
<GID>272</GID>
<name>N_in1</name></connection>
<intersection>366.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-136.5,-94,-87.5,-94</points>
<intersection>-136.5 5</intersection>
<intersection>-87.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-136.5,-94,-136.5,-86.5</points>
<connection>
<GID>238</GID>
<name>OUT_3</name></connection>
<intersection>-94 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-87.5,-94,-87.5,-85.5</points>
<connection>
<GID>240</GID>
<name>IN_3</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-94,-87.5,-84.5</points>
<connection>
<GID>240</GID>
<name>IN_2</name></connection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-136.5,-94,-87.5,-94</points>
<intersection>-136.5 3</intersection>
<intersection>-87.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-136.5,-94,-136.5,-88.5</points>
<connection>
<GID>238</GID>
<name>OUT_2</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362,-11.5,362,-4</points>
<connection>
<GID>281</GID>
<name>OUT</name></connection>
<intersection>-11.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>353,-11.5,362,-11.5</points>
<connection>
<GID>282</GID>
<name>IN_B_0</name></connection>
<intersection>362 0</intersection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-11.5,352,-7.5</points>
<connection>
<GID>282</GID>
<name>IN_B_1</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>358,-7.5,358,-4</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>352,-7.5,358,-7.5</points>
<intersection>352 0</intersection>
<intersection>358 1</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351,-11.5,351,-4</points>
<connection>
<GID>282</GID>
<name>IN_B_2</name></connection>
<intersection>-4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>351,-4,354,-4</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<intersection>351 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-11.5,350,-4</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<connection>
<GID>282</GID>
<name>IN_B_3</name></connection></vsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520.5,-13,520.5,-7.5</points>
<intersection>-13 3</intersection>
<intersection>-7.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>520.5,-13,528,-13</points>
<connection>
<GID>410</GID>
<name>IN_1</name></connection>
<intersection>520.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>513.5,-7.5,520.5,-7.5</points>
<connection>
<GID>325</GID>
<name>OUT_3</name></connection>
<intersection>520.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347.5,-22,347.5,-19.5</points>
<connection>
<GID>282</GID>
<name>OUT_2</name></connection>
<intersection>-22 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>342,-22,347.5,-22</points>
<intersection>342 12</intersection>
<intersection>347.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>342,-25,342,-22</points>
<connection>
<GID>283</GID>
<name>IN_B_2</name></connection>
<intersection>-22 5</intersection></vsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,-23,349.5,-19.5</points>
<connection>
<GID>282</GID>
<name>OUT_0</name></connection>
<intersection>-23 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>344,-23,349.5,-23</points>
<intersection>344 9</intersection>
<intersection>349.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>344,-25,344,-23</points>
<connection>
<GID>283</GID>
<name>IN_B_0</name></connection>
<intersection>-23 5</intersection></vsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341,-25,341,-21.5</points>
<connection>
<GID>283</GID>
<name>IN_B_3</name></connection>
<intersection>-21.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>341,-21.5,346.5,-21.5</points>
<intersection>341 0</intersection>
<intersection>346.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>346.5,-21.5,346.5,-19.5</points>
<connection>
<GID>282</GID>
<name>OUT_3</name></connection>
<intersection>-21.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>348.5,-22.5,348.5,-19.5</points>
<connection>
<GID>282</GID>
<name>OUT_1</name></connection>
<intersection>-22.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>343,-22.5,348.5,-22.5</points>
<intersection>343 6</intersection>
<intersection>348.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>343,-25,343,-22.5</points>
<connection>
<GID>283</GID>
<name>IN_B_1</name></connection>
<intersection>-22.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-94,-87.5,-83.5</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-136.5,-94,-87.5,-94</points>
<intersection>-136.5 3</intersection>
<intersection>-87.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-136.5,-94,-136.5,-90.5</points>
<connection>
<GID>238</GID>
<name>OUT_1</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-94,-87.5,-82.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-136.5,-94,-87.5,-94</points>
<intersection>-136.5 3</intersection>
<intersection>-87.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-136.5,-94,-136.5,-92.5</points>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349,2,349,13.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>13.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>349,13.5,384,13.5</points>
<intersection>349 0</intersection>
<intersection>384 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>384,13.5,384,27.5</points>
<intersection>13.5 2</intersection>
<intersection>27.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>381.5,27.5,384,27.5</points>
<connection>
<GID>246</GID>
<name>OUT_3</name></connection>
<intersection>384 3</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>353,12.5,383.5,12.5</points>
<intersection>353 4</intersection>
<intersection>383.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383.5,12.5,383.5,25.5</points>
<intersection>12.5 1</intersection>
<intersection>25.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>381.5,25.5,383.5,25.5</points>
<connection>
<GID>246</GID>
<name>OUT_2</name></connection>
<intersection>383.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>353,2,353,12.5</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,2,357,11.5</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,11.5,383,11.5</points>
<intersection>357 0</intersection>
<intersection>383 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383,11.5,383,23.5</points>
<intersection>11.5 1</intersection>
<intersection>23.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>381.5,23.5,383,23.5</points>
<connection>
<GID>246</GID>
<name>OUT_1</name></connection>
<intersection>383 2</intersection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361,2,361,10.5</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361,10.5,381.5,10.5</points>
<intersection>361 0</intersection>
<intersection>381.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>381.5,10.5,381.5,21.5</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380.5,2,380.5,9</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380.5,9,400.5,9</points>
<intersection>380.5 0</intersection>
<intersection>400.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>400.5,9,400.5,27</points>
<intersection>9 1</intersection>
<intersection>27 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>396,27,400.5,27</points>
<connection>
<GID>248</GID>
<name>OUT_3</name></connection>
<intersection>400.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384.5,2,384.5,8.5</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384.5,8.5,399.5,8.5</points>
<intersection>384.5 0</intersection>
<intersection>399.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>399.5,8.5,399.5,25</points>
<intersection>8.5 1</intersection>
<intersection>25 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>396,25,399.5,25</points>
<connection>
<GID>248</GID>
<name>OUT_2</name></connection>
<intersection>399.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>388.5,2,388.5,7.5</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>388.5,7.5,398.5,7.5</points>
<intersection>388.5 0</intersection>
<intersection>398.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>398.5,7.5,398.5,23</points>
<intersection>7.5 1</intersection>
<intersection>23 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>396,23,398.5,23</points>
<connection>
<GID>248</GID>
<name>OUT_1</name></connection>
<intersection>398.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>392.5,2,392.5,7</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>392.5,7,397.5,7</points>
<intersection>392.5 0</intersection>
<intersection>397.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>397.5,7,397.5,21</points>
<intersection>7 1</intersection>
<intersection>21 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>396,21,397.5,21</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>397.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361.5,15.5,361.5,27.5</points>
<intersection>15.5 2</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360.5,27.5,361.5,27.5</points>
<connection>
<GID>245</GID>
<name>OUT_3</name></connection>
<intersection>361.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>361.5,15.5,365.5,15.5</points>
<intersection>361.5 0</intersection>
<intersection>365.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>365.5,-25,365.5,15.5</points>
<connection>
<GID>241</GID>
<name>IN_3</name></connection>
<intersection>15.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,-25,366.5,16</points>
<connection>
<GID>241</GID>
<name>IN_2</name></connection>
<intersection>16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>362.5,16,366.5,16</points>
<intersection>362.5 2</intersection>
<intersection>366.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>362.5,16,362.5,25.5</points>
<intersection>16 1</intersection>
<intersection>25.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>360.5,25.5,362.5,25.5</points>
<connection>
<GID>245</GID>
<name>OUT_2</name></connection>
<intersection>362.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363,16.5,363,23.5</points>
<intersection>16.5 2</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360.5,23.5,363,23.5</points>
<connection>
<GID>245</GID>
<name>OUT_1</name></connection>
<intersection>363 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>363,16.5,367.5,16.5</points>
<intersection>363 0</intersection>
<intersection>367.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>367.5,-25,367.5,16.5</points>
<connection>
<GID>241</GID>
<name>IN_1</name></connection>
<intersection>16.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363.5,17,363.5,21.5</points>
<intersection>17 2</intersection>
<intersection>21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360.5,21.5,363.5,21.5</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>363.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>363.5,17,368.5,17</points>
<intersection>363.5 0</intersection>
<intersection>368.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>368.5,-25,368.5,17</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>17 2</intersection></vsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,-25,334,17</points>
<connection>
<GID>283</GID>
<name>IN_3</name></connection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>334,17,350.5,17</points>
<intersection>334 0</intersection>
<intersection>350.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350.5,17,350.5,27.5</points>
<intersection>17 1</intersection>
<intersection>27.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>349,27.5,350.5,27.5</points>
<connection>
<GID>244</GID>
<name>OUT_3</name></connection>
<intersection>350.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335,-25,335,16.5</points>
<connection>
<GID>283</GID>
<name>IN_2</name></connection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>335,16.5,350,16.5</points>
<intersection>335 0</intersection>
<intersection>350 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350,16.5,350,25.5</points>
<intersection>16.5 1</intersection>
<intersection>25.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>349,25.5,350,25.5</points>
<connection>
<GID>244</GID>
<name>OUT_2</name></connection>
<intersection>350 2</intersection></hsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336,-25,336,16</points>
<connection>
<GID>283</GID>
<name>IN_1</name></connection>
<intersection>16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>336,16,349.5,16</points>
<intersection>336 0</intersection>
<intersection>349.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>349.5,16,349.5,23.5</points>
<intersection>16 1</intersection>
<intersection>23.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>349,23.5,349.5,23.5</points>
<connection>
<GID>244</GID>
<name>OUT_1</name></connection>
<intersection>349.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-25,337,15.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>337,15.5,349,15.5</points>
<intersection>337 0</intersection>
<intersection>349 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>349,15.5,349,21.5</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362.5,-40.5,362.5,-35</points>
<connection>
<GID>284</GID>
<name>IN_B_2</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>362.5,-35,370,-35</points>
<intersection>362.5 0</intersection>
<intersection>370 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>370,-49,370,-33</points>
<connection>
<GID>241</GID>
<name>OUT_2</name></connection>
<connection>
<GID>288</GID>
<name>IN_B_2</name></connection>
<intersection>-35 1</intersection></vsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363.5,-40.5,363.5,-36</points>
<connection>
<GID>284</GID>
<name>IN_B_1</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>363.5,-36,371,-36</points>
<intersection>363.5 0</intersection>
<intersection>371 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>371,-49,371,-33</points>
<connection>
<GID>241</GID>
<name>OUT_1</name></connection>
<connection>
<GID>288</GID>
<name>IN_B_1</name></connection>
<intersection>-36 1</intersection></vsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-49,372,-33</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<connection>
<GID>288</GID>
<name>IN_B_0</name></connection>
<intersection>-36.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>364.5,-36.5,372,-36.5</points>
<intersection>364.5 6</intersection>
<intersection>372 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>364.5,-40.5,364.5,-36.5</points>
<connection>
<GID>284</GID>
<name>IN_B_0</name></connection>
<intersection>-36.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361.5,-40.5,361.5,-34.5</points>
<connection>
<GID>284</GID>
<name>IN_B_3</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361.5,-34.5,369,-34.5</points>
<intersection>361.5 0</intersection>
<intersection>369 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>369,-49,369,-33</points>
<connection>
<GID>241</GID>
<name>OUT_3</name></connection>
<connection>
<GID>288</GID>
<name>IN_B_3</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-54.5,-87.5,-42.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-137,-54.5,-87.5,-54.5</points>
<intersection>-137 3</intersection>
<intersection>-87.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-137,-54.5,-137,-51.5</points>
<intersection>-54.5 2</intersection>
<intersection>-51.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-137.5,-51.5,-137,-51.5</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>-137 3</intersection></hsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354.5,-40.5,354.5,-40.5</points>
<connection>
<GID>284</GID>
<name>IN_3</name></connection>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357.5,-40.5,357.5,-40.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-53,-87.5,-43.5</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-137,-53,-87.5,-53</points>
<intersection>-137 3</intersection>
<intersection>-87.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-137,-53,-137,-49.5</points>
<intersection>-53 2</intersection>
<intersection>-49.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-137.5,-49.5,-137,-49.5</points>
<connection>
<GID>232</GID>
<name>OUT_1</name></connection>
<intersection>-137 3</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331,-40,331,-34.5</points>
<connection>
<GID>290</GID>
<name>IN_B_2</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>331,-34.5,338.5,-34.5</points>
<intersection>331 0</intersection>
<intersection>338.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>338.5,-49,338.5,-33</points>
<connection>
<GID>283</GID>
<name>OUT_2</name></connection>
<connection>
<GID>297</GID>
<name>IN_B_2</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,-40,332,-35.5</points>
<connection>
<GID>290</GID>
<name>IN_B_1</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>332,-35.5,339.5,-35.5</points>
<intersection>332 0</intersection>
<intersection>339.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>339.5,-49,339.5,-33</points>
<connection>
<GID>283</GID>
<name>OUT_1</name></connection>
<connection>
<GID>297</GID>
<name>IN_B_1</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>340.5,-49,340.5,-33</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<connection>
<GID>297</GID>
<name>IN_B_0</name></connection>
<intersection>-36 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>333,-36,340.5,-36</points>
<intersection>333 6</intersection>
<intersection>340.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>333,-40,333,-36</points>
<connection>
<GID>290</GID>
<name>IN_B_0</name></connection>
<intersection>-36 4</intersection></vsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,-40,330,-34</points>
<connection>
<GID>290</GID>
<name>IN_B_3</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>330,-34,337.5,-34</points>
<intersection>330 0</intersection>
<intersection>337.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>337.5,-49,337.5,-33</points>
<connection>
<GID>283</GID>
<name>OUT_3</name></connection>
<connection>
<GID>297</GID>
<name>IN_B_3</name></connection>
<intersection>-34 1</intersection></vsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323,-40,323,-40</points>
<connection>
<GID>290</GID>
<name>IN_3</name></connection>
<connection>
<GID>295</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520.5,-9,520.5,-6.5</points>
<intersection>-9 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,-6.5,520.5,-6.5</points>
<connection>
<GID>325</GID>
<name>OUT_2</name></connection>
<intersection>520.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>520.5,-9,528,-9</points>
<connection>
<GID>409</GID>
<name>IN_1</name></connection>
<intersection>520.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520.5,-5.5,520.5,-5</points>
<intersection>-5.5 1</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,-5.5,520.5,-5.5</points>
<connection>
<GID>325</GID>
<name>OUT_1</name></connection>
<intersection>520.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>520.5,-5,528,-5</points>
<connection>
<GID>408</GID>
<name>IN_1</name></connection>
<intersection>520.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>314.5,-48,332.5,-48</points>
<intersection>314.5 8</intersection>
<intersection>320 3</intersection>
<intersection>331.5 13</intersection>
<intersection>332.5 14</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>320,-48,320,-46</points>
<connection>
<GID>290</GID>
<name>A_less_B</name></connection>
<intersection>-48 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>314.5,-52.5,314.5,-48</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>-48 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>331.5,-49,331.5,-48</points>
<connection>
<GID>297</GID>
<name>IN_2</name></connection>
<intersection>-48 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>332.5,-49,332.5,-48</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>-48 1</intersection></vsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>349,-58.5,372.5,-58.5</points>
<connection>
<GID>307</GID>
<name>OUT_0</name></connection>
<intersection>349 26</intersection>
<intersection>360.5 39</intersection>
<intersection>364.5 27</intersection>
<intersection>368.5 28</intersection>
<intersection>372.5 29</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>349,-69,349,-58.5</points>
<intersection>-69 30</intersection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>364.5,-60,364.5,-58.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>368.5,-60,368.5,-58.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>372.5,-60,372.5,-58.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>349,-69,357.5,-69</points>
<intersection>349 26</intersection>
<intersection>355.5 42</intersection>
<intersection>357.5 32</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>357.5,-70,357.5,-69</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>-69 30</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>360.5,-60,360.5,-58.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>355.5,-70,355.5,-69</points>
<connection>
<GID>302</GID>
<name>IN_3</name></connection>
<intersection>-69 30</intersection></vsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,-74.5,-51,-74.5</points>
<connection>
<GID>275</GID>
<name>IN_B_0</name></connection>
<intersection>-79 9</intersection>
<intersection>-72.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-72.5,-74.5,-72.5,-59.5</points>
<intersection>-74.5 1</intersection>
<intersection>-59.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-72.5,-59.5,-28.5,-59.5</points>
<connection>
<GID>273</GID>
<name>IN_B_0</name></connection>
<intersection>-72.5 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-79,-79,-79,-74.5</points>
<intersection>-79 12</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-79.5,-79,-79,-79</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<intersection>-79 9</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,-76.5,-51,-76.5</points>
<connection>
<GID>275</GID>
<name>IN_B_2</name></connection>
<intersection>-76.5 8</intersection>
<intersection>-70.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-70.5,-76.5,-70.5,-61.5</points>
<intersection>-76.5 1</intersection>
<intersection>-61.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-70.5,-61.5,-28.5,-61.5</points>
<connection>
<GID>273</GID>
<name>IN_B_2</name></connection>
<intersection>-70.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-76.5,-81,-76.5,-76.5</points>
<intersection>-81 9</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-79.5,-81,-76.5,-81</points>
<connection>
<GID>240</GID>
<name>OUT_2</name></connection>
<intersection>-76.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-77.5,-75.5,-51,-75.5</points>
<connection>
<GID>275</GID>
<name>IN_B_1</name></connection>
<intersection>-77.5 10</intersection>
<intersection>-71.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-71.5,-75.5,-71.5,-60.5</points>
<intersection>-75.5 1</intersection>
<intersection>-60.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-71.5,-60.5,-28.5,-60.5</points>
<connection>
<GID>273</GID>
<name>IN_B_1</name></connection>
<intersection>-71.5 8</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-77.5,-80,-77.5,-75.5</points>
<intersection>-80 14</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-79.5,-80,-77.5,-80</points>
<connection>
<GID>240</GID>
<name>OUT_1</name></connection>
<intersection>-77.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>347,-28,362.5,-28</points>
<connection>
<GID>241</GID>
<name>carry_out</name></connection>
<connection>
<GID>283</GID>
<name>carry_in</name></connection>
<intersection>348 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>348,-46.5,348,-28</points>
<connection>
<GID>400</GID>
<name>IN_1</name></connection>
<intersection>-28 1</intersection></vsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353.5,-67.5,353.5,-48</points>
<intersection>-67.5 1</intersection>
<intersection>-54.5 14</intersection>
<intersection>-48 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353.5,-67.5,370,-67.5</points>
<intersection>353.5 0</intersection>
<intersection>370 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>370,-73,370,-67.5</points>
<intersection>-73 3</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>368.5,-73,370,-73</points>
<connection>
<GID>302</GID>
<name>carry_in</name></connection>
<intersection>370 2</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>353.5,-48,364,-48</points>
<intersection>353.5 0</intersection>
<intersection>363 12</intersection>
<intersection>364 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>364,-49,364,-48</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<intersection>-48 8</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>363,-49,363,-48</points>
<connection>
<GID>288</GID>
<name>IN_2</name></connection>
<intersection>-48 8</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>349,-54.5,353.5,-54.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>349 18</intersection>
<intersection>353.5 0</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>349,-54.5,349,-52.5</points>
<connection>
<GID>400</GID>
<name>OUT</name></connection>
<intersection>-54.5 14</intersection></vsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>368,-69,368,-66.5</points>
<intersection>-69 3</intersection>
<intersection>-66.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>371.5,-66.5,371.5,-66</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>368,-66.5,371.5,-66.5</points>
<intersection>368 0</intersection>
<intersection>371.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>365.5,-69,368,-69</points>
<intersection>365.5 4</intersection>
<intersection>368 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>365.5,-70,365.5,-69</points>
<connection>
<GID>302</GID>
<name>IN_B_0</name></connection>
<intersection>-69 3</intersection></vsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>364.5,-70,364.5,-68.5</points>
<connection>
<GID>302</GID>
<name>IN_B_1</name></connection>
<intersection>-68.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>367.5,-68.5,367.5,-66</points>
<connection>
<GID>300</GID>
<name>OUT</name></connection>
<intersection>-68.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>364.5,-68.5,367.5,-68.5</points>
<intersection>364.5 0</intersection>
<intersection>367.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363.5,-70,363.5,-66</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<connection>
<GID>302</GID>
<name>IN_B_2</name></connection></vsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361,-69,361,-66</points>
<intersection>-69 3</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>359.5,-66,361,-66</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<intersection>361 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>361,-69,362.5,-69</points>
<intersection>361 0</intersection>
<intersection>362.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>362.5,-70,362.5,-69</points>
<connection>
<GID>302</GID>
<name>IN_B_3</name></connection>
<intersection>-69 3</intersection></vsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-74,-77.5,-51,-77.5</points>
<connection>
<GID>275</GID>
<name>IN_B_3</name></connection>
<intersection>-74 8</intersection>
<intersection>-69 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-69,-77.5,-69,-62.5</points>
<intersection>-77.5 1</intersection>
<intersection>-62.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-69,-62.5,-28.5,-62.5</points>
<connection>
<GID>273</GID>
<name>IN_B_3</name></connection>
<intersection>-69 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-74,-82,-74,-77.5</points>
<intersection>-82 9</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-79.5,-82,-74,-82</points>
<connection>
<GID>240</GID>
<name>OUT_3</name></connection>
<intersection>-74 8</intersection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>358.5,-60,358.5,-57</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>358.5,-57,365.5,-57</points>
<connection>
<GID>288</GID>
<name>OUT_3</name></connection>
<intersection>358.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,-57.5,366.5,-57</points>
<connection>
<GID>288</GID>
<name>OUT_2</name></connection>
<intersection>-57.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>362.5,-60,362.5,-57.5</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>362.5,-57.5,366.5,-57.5</points>
<intersection>362.5 1</intersection>
<intersection>366.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,-60,366.5,-58</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>367.5,-58,367.5,-57</points>
<connection>
<GID>288</GID>
<name>OUT_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>366.5,-58,367.5,-58</points>
<intersection>366.5 0</intersection>
<intersection>367.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370.5,-60,370.5,-58</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>368.5,-58,368.5,-57</points>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>368.5,-58,370.5,-58</points>
<intersection>368.5 1</intersection>
<intersection>370.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520.5,-4.5,520.5,-1</points>
<intersection>-4.5 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,-4.5,520.5,-4.5</points>
<connection>
<GID>325</GID>
<name>OUT_0</name></connection>
<intersection>520.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>520.5,-1,528,-1</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<intersection>520.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>513.5,8.5,528,8.5</points>
<connection>
<GID>406</GID>
<name>IN_1</name></connection>
<connection>
<GID>313</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>521,9.5,521,13</points>
<intersection>9.5 1</intersection>
<intersection>13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,9.5,521,9.5</points>
<connection>
<GID>313</GID>
<name>OUT_2</name></connection>
<intersection>521 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>521,13,528,13</points>
<connection>
<GID>405</GID>
<name>IN_1</name></connection>
<intersection>521 0</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>519.5,10.5,519.5,18.5</points>
<intersection>10.5 1</intersection>
<intersection>18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,10.5,519.5,10.5</points>
<connection>
<GID>313</GID>
<name>OUT_1</name></connection>
<intersection>519.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>519.5,18.5,528,18.5</points>
<connection>
<GID>404</GID>
<name>IN_1</name></connection>
<intersection>519.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520,11.5,520,29.5</points>
<intersection>11.5 1</intersection>
<intersection>29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,11.5,520,11.5</points>
<connection>
<GID>313</GID>
<name>OUT_0</name></connection>
<intersection>520 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>520,29.5,528,29.5</points>
<connection>
<GID>403</GID>
<name>IN_1</name></connection>
<intersection>520 0</intersection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509.5,20.5,509.5,22</points>
<connection>
<GID>312</GID>
<name>carry_out</name></connection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>509.5,20.5,528,20.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>509.5 0</intersection>
<intersection>525 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>525,-11,525,31.5</points>
<intersection>-11 33</intersection>
<intersection>-7 31</intersection>
<intersection>-3 30</intersection>
<intersection>1 29</intersection>
<intersection>10.5 3</intersection>
<intersection>15 6</intersection>
<intersection>20.5 1</intersection>
<intersection>31.5 28</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>525,10.5,528,10.5</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>525,15,528,15</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>525,31.5,528,31.5</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>525,1,528,1</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>525,-3,528,-3</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>525,-7,528,-7</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>525,-11,528,-11</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>534,30.5,545.5,30.5</points>
<connection>
<GID>403</GID>
<name>OUT</name></connection>
<connection>
<GID>411</GID>
<name>IN_B_0</name></connection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51,-84.5,-51,-84.5</points>
<connection>
<GID>275</GID>
<name>IN_3</name></connection>
<connection>
<GID>285</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88,-52,-88,-44.5</points>
<intersection>-52 1</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-137,-52,-88,-52</points>
<intersection>-137 3</intersection>
<intersection>-88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-88,-44.5,-87.5,-44.5</points>
<connection>
<GID>236</GID>
<name>IN_2</name></connection>
<intersection>-88 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-137,-52,-137,-47.5</points>
<intersection>-52 1</intersection>
<intersection>-47.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-137.5,-47.5,-137,-47.5</points>
<connection>
<GID>232</GID>
<name>OUT_2</name></connection>
<intersection>-137 3</intersection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-137,-51,-87.5,-51</points>
<intersection>-137 3</intersection>
<intersection>-87.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-87.5,-51,-87.5,-45.5</points>
<connection>
<GID>236</GID>
<name>IN_3</name></connection>
<intersection>-51 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>-137,-51,-137,-45.5</points>
<intersection>-51 1</intersection>
<intersection>-45.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-137.5,-45.5,-137,-45.5</points>
<connection>
<GID>232</GID>
<name>OUT_3</name></connection>
<intersection>-137 3</intersection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-1,-77,-1,-77</points>
<connection>
<GID>304</GID>
<name>N_in2</name></connection>
<connection>
<GID>317</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-1,-79,-1,-79</points>
<connection>
<GID>317</GID>
<name>N_in2</name></connection>
<connection>
<GID>318</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>537.5,19.5,537.5,29.5</points>
<intersection>19.5 2</intersection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>537.5,29.5,545.5,29.5</points>
<connection>
<GID>411</GID>
<name>IN_B_1</name></connection>
<intersection>537.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>534,19.5,537.5,19.5</points>
<connection>
<GID>404</GID>
<name>OUT</name></connection>
<intersection>537.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84.5,-72.5,-84.5,-48.5</points>
<connection>
<GID>240</GID>
<name>carry_in</name></connection>
<connection>
<GID>236</GID>
<name>carry_out</name></connection>
<intersection>-55 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-84.5,-55,-75.5,-55</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<intersection>-84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-29,-5.5,-26</points>
<connection>
<GID>305</GID>
<name>IN_3</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-29,-5.5,-29</points>
<connection>
<GID>242</GID>
<name>OUT_3</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-28,-5.5,-27</points>
<connection>
<GID>305</GID>
<name>IN_2</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-28,-5.5,-28</points>
<connection>
<GID>242</GID>
<name>OUT_2</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-5.5,-28,-5.5,-27</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>-27 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-20.5,-27,-5.5,-27</points>
<connection>
<GID>242</GID>
<name>OUT_1</name></connection>
<intersection>-5.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-29,-5.5,-26</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-26,-5.5,-26</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-48.5,-52.5,-46,-52.5</points>
<intersection>-48.5 6</intersection>
<intersection>-46 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-48.5,-52.5,-48.5,-52</points>
<connection>
<GID>252</GID>
<name>A_less_B</name></connection>
<intersection>-52.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-46,-52.5,-46,-52</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>-52.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-66,-4,-63</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-63,-4,-63</points>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-65,-21,-64</points>
<intersection>-65 1</intersection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-65,-4,-65</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-64,-20.5,-64</points>
<connection>
<GID>273</GID>
<name>OUT_1</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-65,-4,-64</points>
<connection>
<GID>309</GID>
<name>IN_2</name></connection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-65,-4,-65</points>
<connection>
<GID>273</GID>
<name>OUT_2</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-66,-3.5,-63</points>
<intersection>-66 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-66,-3.5,-66</points>
<connection>
<GID>273</GID>
<name>OUT_3</name></connection>
<intersection>-3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-63,-3.5,-63</points>
<connection>
<GID>309</GID>
<name>IN_3</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45,-90,-45,-87.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<connection>
<GID>275</GID>
<name>A_less_B</name></connection></vsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-81,-1,-81</points>
<connection>
<GID>319</GID>
<name>N_in3</name></connection>
<connection>
<GID>318</GID>
<name>N_in2</name></connection>
<intersection>-1.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1.5,-81,-1.5,-80</points>
<intersection>-81 1</intersection>
<intersection>-80 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-2,-80,-1.5,-80</points>
<connection>
<GID>318</GID>
<name>N_in0</name></connection>
<intersection>-1.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,-56.5,-25.5,-35.5</points>
<connection>
<GID>273</GID>
<name>carry_in</name></connection>
<connection>
<GID>242</GID>
<name>carry_out</name></connection>
<intersection>-55.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-63.5,-55.5,-25.5,-55.5</points>
<intersection>-63.5 9</intersection>
<intersection>-25.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-63.5,-82.5,-63.5,-55.5</points>
<intersection>-82.5 10</intersection>
<intersection>-55.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-63.5,-82.5,-58.5,-82.5</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>-63.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-58.5,-80.5,-58.5,-80.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>316</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-52.5,-81.5,-51,-81.5</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<connection>
<GID>275</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-75,4.5,-11</points>
<intersection>-75 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-82.5,-11,4.5,-11</points>
<connection>
<GID>320</GID>
<name>OUT</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,-75,4.5,-75</points>
<connection>
<GID>304</GID>
<name>N_in3</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45,-46,-45,-33.5</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>-37.5 21</intersection>
<intersection>-33.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-45,-33.5,-36,-33.5</points>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<intersection>-45 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-45,-37.5,-36,-37.5</points>
<connection>
<GID>323</GID>
<name>IN_1</name></connection>
<intersection>-45 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-36.5,-29,-31.5</points>
<intersection>-36.5 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,-31.5,-28.5,-31.5</points>
<connection>
<GID>242</GID>
<name>IN_2</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-30,-36.5,-29,-36.5</points>
<connection>
<GID>323</GID>
<name>OUT</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-32.5,-29.5,-30.5</points>
<intersection>-32.5 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-30.5,-28.5,-30.5</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-30,-32.5,-29.5,-32.5</points>
<connection>
<GID>322</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-29.5,-29.5,-28.5</points>
<intersection>-29.5 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-29.5,-28.5,-29.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-30,-28.5,-29.5,-28.5</points>
<connection>
<GID>321</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-40.5,-28.5,-32.5</points>
<connection>
<GID>242</GID>
<name>IN_3</name></connection>
<intersection>-40.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-30,-40.5,-28.5,-40.5</points>
<connection>
<GID>324</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>538.5,14,538.5,28.5</points>
<intersection>14 1</intersection>
<intersection>28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534,14,538.5,14</points>
<connection>
<GID>405</GID>
<name>OUT</name></connection>
<intersection>538.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>538.5,28.5,545.5,28.5</points>
<connection>
<GID>411</GID>
<name>IN_B_2</name></connection>
<intersection>538.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-29.5,-36,-29.5</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<connection>
<GID>321</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-41.5,-36,-41.5</points>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<connection>
<GID>324</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-81.5,-38,-69.5</points>
<intersection>-81.5 28</intersection>
<intersection>-73.5 21</intersection>
<intersection>-69.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-38,-69.5,-35.5,-69.5</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>-38 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-38,-73.5,-35.5,-73.5</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<intersection>-38 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-38,-81.5,-36,-81.5</points>
<connection>
<GID>329</GID>
<name>OUT</name></connection>
<intersection>-38 0</intersection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-65.5,-35.5,-65.5</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<connection>
<GID>229</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-77.5,-35.5,-77.5</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<connection>
<GID>234</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539.5,9.5,539.5,27.5</points>
<intersection>9.5 2</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>539.5,27.5,545.5,27.5</points>
<connection>
<GID>411</GID>
<name>IN_B_3</name></connection>
<intersection>539.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>534,9.5,539.5,9.5</points>
<connection>
<GID>406</GID>
<name>OUT</name></connection>
<intersection>539.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-105.5,-77.5,-105.5,-16.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<connection>
<GID>271</GID>
<name>OUT</name></connection>
<intersection>-36.5 101</intersection>
<intersection>-32.5 39</intersection>
<intersection>-28.5 29</intersection>
<intersection>-24.5 28</intersection>
<intersection>-16.5 30</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-105.5,-24.5,-104.5,-24.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-105.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-105.5,-28.5,-104.5,-28.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-105.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-105.5,-16.5,-25.5,-16.5</points>
<intersection>-105.5 0</intersection>
<intersection>-84.5 233</intersection>
<intersection>-40 37</intersection>
<intersection>-25.5 226</intersection></hsegment>
<vsegment>
<ID>37</ID>
<points>-40,-88,-40,-16.5</points>
<intersection>-88 240</intersection>
<intersection>-75.5 90</intersection>
<intersection>-71.5 98</intersection>
<intersection>-67.5 95</intersection>
<intersection>-63.5 96</intersection>
<intersection>-39.5 237</intersection>
<intersection>-35.5 48</intersection>
<intersection>-31.5 45</intersection>
<intersection>-27.5 228</intersection>
<intersection>-16.5 30</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>-105.5,-32.5,-104.5,-32.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>-105.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>-40,-31.5,-36,-31.5</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-40,-35.5,-36,-35.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>90</ID>
<points>-40,-75.5,-35.5,-75.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>95</ID>
<points>-40,-67.5,-35.5,-67.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>96</ID>
<points>-40,-63.5,-35.5,-63.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>98</ID>
<points>-40,-71.5,-35.5,-71.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>101</ID>
<points>-105.5,-36.5,-104.5,-36.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>-105.5 0</intersection></hsegment>
<vsegment>
<ID>226</ID>
<points>-25.5,-19.5,-25.5,-16.5</points>
<connection>
<GID>242</GID>
<name>carry_in</name></connection>
<intersection>-16.5 30</intersection></vsegment>
<hsegment>
<ID>228</ID>
<points>-40,-27.5,-36,-27.5</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<vsegment>
<ID>233</ID>
<points>-84.5,-53,-84.5,-16.5</points>
<connection>
<GID>236</GID>
<name>carry_in</name></connection>
<intersection>-53 234</intersection>
<intersection>-16.5 30</intersection></vsegment>
<hsegment>
<ID>234</ID>
<points>-84.5,-53,-75.5,-53</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>-84.5 233</intersection></hsegment>
<hsegment>
<ID>237</ID>
<points>-40,-39.5,-36,-39.5</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>240</ID>
<points>-40,-88,-37,-88</points>
<intersection>-40 37</intersection>
<intersection>-37 241</intersection></hsegment>
<vsegment>
<ID>241</ID>
<points>-37,-88,-37,-87.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>-88 240</intersection></vsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>537,0,537,8.5</points>
<intersection>0 1</intersection>
<intersection>8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534,0,537,0</points>
<connection>
<GID>407</GID>
<name>OUT</name></connection>
<intersection>537 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>537,8.5,545.5,8.5</points>
<connection>
<GID>412</GID>
<name>IN_B_0</name></connection>
<intersection>537 0</intersection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>536,-4,536,7.5</points>
<intersection>-4 1</intersection>
<intersection>7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534,-4,536,-4</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>536 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>536,7.5,545.5,7.5</points>
<connection>
<GID>412</GID>
<name>IN_B_1</name></connection>
<intersection>536 0</intersection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>538,-8,538,6.5</points>
<intersection>-8 1</intersection>
<intersection>6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534,-8,538,-8</points>
<connection>
<GID>409</GID>
<name>OUT</name></connection>
<intersection>538 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>538,6.5,545.5,6.5</points>
<connection>
<GID>412</GID>
<name>IN_B_2</name></connection>
<intersection>538 0</intersection></hsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-76.5,-28.5,-69.5</points>
<connection>
<GID>273</GID>
<name>IN_3</name></connection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,-76.5,-28.5,-76.5</points>
<connection>
<GID>234</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539.5,-12,539.5,5.5</points>
<intersection>-12 3</intersection>
<intersection>5.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>534,-12,539.5,-12</points>
<connection>
<GID>410</GID>
<name>OUT</name></connection>
<intersection>539.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>539.5,5.5,545.5,5.5</points>
<connection>
<GID>412</GID>
<name>IN_B_3</name></connection>
<intersection>539.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-66.5,-29,-64.5</points>
<intersection>-66.5 1</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,-66.5,-28.5,-66.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,-64.5,-29,-64.5</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-68.5,-29.5,-67.5</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-67.5,-28.5,-67.5</points>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>538,-14.5,545.5,-14.5</points>
<intersection>538 3</intersection>
<intersection>545.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>538,-18,538,-14.5</points>
<connection>
<GID>311</GID>
<name>OUT_7</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>545.5,-14.5,545.5,-1.5</points>
<connection>
<GID>412</GID>
<name>IN_3</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-38.5,-106.5,-32</points>
<intersection>-38.5 5</intersection>
<intersection>-32 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-110.5,-32,-106.5,-32</points>
<connection>
<GID>227</GID>
<name>OUT_3</name></connection>
<intersection>-106.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106.5,-38.5,-104.5,-38.5</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-34.5,-106.5,-34</points>
<intersection>-34.5 5</intersection>
<intersection>-34 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-110.5,-34,-106.5,-34</points>
<connection>
<GID>227</GID>
<name>OUT_2</name></connection>
<intersection>-106.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106.5,-34.5,-104.5,-34.5</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-36,-106.5,-30.5</points>
<intersection>-36 4</intersection>
<intersection>-30.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-110.5,-36,-106.5,-36</points>
<connection>
<GID>227</GID>
<name>OUT_1</name></connection>
<intersection>-106.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106.5,-30.5,-104.5,-30.5</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-38,-106.5,-26.5</points>
<intersection>-38 4</intersection>
<intersection>-26.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-110.5,-38,-106.5,-38</points>
<connection>
<GID>227</GID>
<name>OUT_0</name></connection>
<intersection>-106.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106.5,-26.5,-104.5,-26.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>541.5,-19,541.5,-0.5</points>
<intersection>-19 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-19,541.5,-19</points>
<connection>
<GID>311</GID>
<name>OUT_6</name></connection>
<intersection>541.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>541.5,-0.5,545.5,-0.5</points>
<connection>
<GID>412</GID>
<name>IN_2</name></connection>
<intersection>541.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>542,-20,542,0.5</points>
<intersection>-20 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-20,542,-20</points>
<connection>
<GID>311</GID>
<name>OUT_5</name></connection>
<intersection>542 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>542,0.5,545.5,0.5</points>
<connection>
<GID>412</GID>
<name>IN_1</name></connection>
<intersection>542 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-21,540.5,1.5</points>
<intersection>-21 1</intersection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-21,540.5,-21</points>
<connection>
<GID>311</GID>
<name>OUT_4</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,1.5,545.5,1.5</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>540.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>544.5,-22,544.5,20.5</points>
<intersection>-22 1</intersection>
<intersection>20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-22,544.5,-22</points>
<connection>
<GID>311</GID>
<name>OUT_3</name></connection>
<intersection>544.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>544.5,20.5,545.5,20.5</points>
<connection>
<GID>411</GID>
<name>IN_3</name></connection>
<intersection>544.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107.5,-79.5,-107.5,-73</points>
<intersection>-79.5 3</intersection>
<intersection>-73 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-107.5,-79.5,-105.5,-79.5</points>
<connection>
<GID>226</GID>
<name>IN_1</name></connection>
<intersection>-107.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-112,-73,-107.5,-73</points>
<connection>
<GID>235</GID>
<name>OUT_3</name></connection>
<intersection>-107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107.5,-75.5,-107.5,-75</points>
<intersection>-75.5 3</intersection>
<intersection>-75 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-107.5,-75.5,-105.5,-75.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>-107.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-112,-75,-107.5,-75</points>
<connection>
<GID>235</GID>
<name>OUT_2</name></connection>
<intersection>-107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107.5,-77,-107.5,-71.5</points>
<intersection>-77 4</intersection>
<intersection>-71.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-107.5,-71.5,-105.5,-71.5</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>-107.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-112,-77,-107.5,-77</points>
<connection>
<GID>235</GID>
<name>OUT_1</name></connection>
<intersection>-107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107.5,-79,-107.5,-67.5</points>
<intersection>-79 4</intersection>
<intersection>-67.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-107.5,-67.5,-105.5,-67.5</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>-107.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-112,-79,-107.5,-79</points>
<connection>
<GID>235</GID>
<name>OUT_0</name></connection>
<intersection>-107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84.5,-92,-84.5,-88.5</points>
<connection>
<GID>240</GID>
<name>carry_out</name></connection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-84.5,-92,-45,-92</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>-84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93,-35.5,-93,-25.5</points>
<intersection>-35.5 1</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93,-35.5,-87.5,-35.5</points>
<connection>
<GID>236</GID>
<name>IN_B_0</name></connection>
<intersection>-93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-98.5,-25.5,-93,-25.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>-93 0</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93,-36.5,-93,-29.5</points>
<intersection>-36.5 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-98.5,-29.5,-93,-29.5</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>-93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-93,-36.5,-87.5,-36.5</points>
<connection>
<GID>236</GID>
<name>IN_B_1</name></connection>
<intersection>-93 0</intersection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93,-37.5,-93,-33.5</points>
<intersection>-37.5 1</intersection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93,-37.5,-87.5,-37.5</points>
<connection>
<GID>236</GID>
<name>IN_B_2</name></connection>
<intersection>-93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-98.5,-33.5,-93,-33.5</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>-93 0</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93,-38.5,-93,-37.5</points>
<intersection>-38.5 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-98.5,-37.5,-93,-37.5</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>-93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-93,-38.5,-87.5,-38.5</points>
<connection>
<GID>236</GID>
<name>IN_B_3</name></connection>
<intersection>-93 0</intersection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93.5,-75.5,-93.5,-66.5</points>
<intersection>-75.5 1</intersection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93.5,-75.5,-87.5,-75.5</points>
<connection>
<GID>240</GID>
<name>IN_B_0</name></connection>
<intersection>-93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-99.5,-66.5,-93.5,-66.5</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>-93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93.5,-76.5,-93.5,-70.5</points>
<intersection>-76.5 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-99.5,-70.5,-93.5,-70.5</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<intersection>-93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-93.5,-76.5,-87.5,-76.5</points>
<connection>
<GID>240</GID>
<name>IN_B_1</name></connection>
<intersection>-93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93.5,-77.5,-93.5,-74.5</points>
<intersection>-77.5 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93.5,-77.5,-87.5,-77.5</points>
<connection>
<GID>240</GID>
<name>IN_B_2</name></connection>
<intersection>-93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-99.5,-74.5,-93.5,-74.5</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<intersection>-93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-99.5,-78.5,-87.5,-78.5</points>
<connection>
<GID>226</GID>
<name>OUT</name></connection>
<connection>
<GID>240</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-54,-44,-52</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,-54,-44,-54</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>543.5,-23,543.5,21.5</points>
<intersection>-23 1</intersection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-23,543.5,-23</points>
<connection>
<GID>311</GID>
<name>OUT_2</name></connection>
<intersection>543.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>543.5,21.5,545.5,21.5</points>
<connection>
<GID>411</GID>
<name>IN_2</name></connection>
<intersection>543.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>542.5,-24,542.5,22.5</points>
<intersection>-24 1</intersection>
<intersection>22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-24,542.5,-24</points>
<connection>
<GID>311</GID>
<name>OUT_1</name></connection>
<intersection>542.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>542.5,22.5,545.5,22.5</points>
<connection>
<GID>411</GID>
<name>IN_1</name></connection>
<intersection>542.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>541,-25,541,23.5</points>
<intersection>-25 1</intersection>
<intersection>23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-25,541,-25</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<intersection>541 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>541,23.5,545.5,23.5</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>541 0</intersection></hsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-91,-35,-87.5</points>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-91,-35,-91</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,-12.5,-268,-12</points>
<connection>
<GID>356</GID>
<name>IN_1</name></connection>
<connection>
<GID>354</GID>
<name>OUT_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-268,-12,-250,-12</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-266,-14,-266,-12.5</points>
<connection>
<GID>337</GID>
<name>OUT_0</name></connection>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-266,-14,-250,-14</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<intersection>-266 0</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-241,-41,-216,-41</points>
<connection>
<GID>343</GID>
<name>OUT_0</name></connection>
<connection>
<GID>350</GID>
<name>IN_B_0</name></connection>
<intersection>-236.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-236.5,-41,-236.5,-24.5</points>
<intersection>-41 1</intersection>
<intersection>-24.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-236.5,-24.5,-190,-24.5</points>
<connection>
<GID>346</GID>
<name>IN_B_0</name></connection>
<intersection>-236.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-241,-43,-216,-43</points>
<connection>
<GID>343</GID>
<name>OUT_2</name></connection>
<connection>
<GID>350</GID>
<name>IN_B_2</name></connection>
<intersection>-234.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-234.5,-43,-234.5,-26.5</points>
<intersection>-43 1</intersection>
<intersection>-26.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-234.5,-26.5,-190,-26.5</points>
<connection>
<GID>346</GID>
<name>IN_B_2</name></connection>
<intersection>-234.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-241,-42,-216,-42</points>
<connection>
<GID>343</GID>
<name>OUT_1</name></connection>
<connection>
<GID>350</GID>
<name>IN_B_1</name></connection>
<intersection>-235.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-235.5,-42,-235.5,-25.5</points>
<intersection>-42 1</intersection>
<intersection>-25.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-235.5,-25.5,-190,-25.5</points>
<connection>
<GID>346</GID>
<name>IN_B_1</name></connection>
<intersection>-235.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-241,-44,-216,-44</points>
<connection>
<GID>343</GID>
<name>OUT_3</name></connection>
<connection>
<GID>350</GID>
<name>IN_B_3</name></connection>
<intersection>-233 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-233,-44,-233,-27.5</points>
<intersection>-44 1</intersection>
<intersection>-27.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-233,-27.5,-190,-27.5</points>
<connection>
<GID>346</GID>
<name>IN_B_3</name></connection>
<intersection>-233 6</intersection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-221,-51,-216,-51</points>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection>
<connection>
<GID>350</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-220.5,-48,-216,-48</points>
<connection>
<GID>352</GID>
<name>OUT_0</name></connection>
<connection>
<GID>350</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-298,-96,-249,-96</points>
<intersection>-298 5</intersection>
<intersection>-249 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-298,-96,-298,-88.5</points>
<connection>
<GID>344</GID>
<name>OUT_3</name></connection>
<intersection>-96 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-249,-96,-249,-87.5</points>
<connection>
<GID>345</GID>
<name>IN_3</name></connection>
<intersection>-96 1</intersection></vsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249,-96,-249,-86.5</points>
<connection>
<GID>345</GID>
<name>IN_2</name></connection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-298,-96,-249,-96</points>
<intersection>-298 3</intersection>
<intersection>-249 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-298,-96,-298,-90.5</points>
<connection>
<GID>344</GID>
<name>OUT_2</name></connection>
<intersection>-96 1</intersection></vsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249,-96,-249,-85.5</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-298,-96,-249,-96</points>
<intersection>-298 3</intersection>
<intersection>-249 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-298,-96,-298,-92.5</points>
<connection>
<GID>344</GID>
<name>OUT_1</name></connection>
<intersection>-96 1</intersection></vsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249,-96,-249,-84.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-298,-96,-249,-96</points>
<intersection>-298 3</intersection>
<intersection>-249 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-298,-96,-298,-94.5</points>
<connection>
<GID>344</GID>
<name>OUT_0</name></connection>
<intersection>-96 1</intersection></vsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249,-56.5,-249,-44.5</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-298.5,-56.5,-249,-56.5</points>
<intersection>-298.5 3</intersection>
<intersection>-249 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-298.5,-57,-298.5,-56.5</points>
<connection>
<GID>339</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249,-55,-249,-45.5</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-298.5,-55,-249,-55</points>
<connection>
<GID>339</GID>
<name>OUT_1</name></connection>
<intersection>-249 0</intersection></hsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-240.5,-76.5,-214,-76.5</points>
<connection>
<GID>359</GID>
<name>IN_B_0</name></connection>
<intersection>-240.5 9</intersection>
<intersection>-234 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-234,-76.5,-234,-61.5</points>
<intersection>-76.5 1</intersection>
<intersection>-61.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-234,-61.5,-190,-61.5</points>
<connection>
<GID>358</GID>
<name>IN_B_0</name></connection>
<intersection>-234 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-240.5,-81,-240.5,-76.5</points>
<intersection>-81 12</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-241,-81,-240.5,-81</points>
<connection>
<GID>345</GID>
<name>OUT_0</name></connection>
<intersection>-240.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-238,-78.5,-214,-78.5</points>
<connection>
<GID>359</GID>
<name>IN_B_2</name></connection>
<intersection>-238 8</intersection>
<intersection>-232 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-232,-78.5,-232,-63.5</points>
<intersection>-78.5 1</intersection>
<intersection>-63.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-232,-63.5,-190,-63.5</points>
<connection>
<GID>358</GID>
<name>IN_B_2</name></connection>
<intersection>-232 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-238,-83,-238,-78.5</points>
<intersection>-83 9</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-241,-83,-238,-83</points>
<connection>
<GID>345</GID>
<name>OUT_2</name></connection>
<intersection>-238 8</intersection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-239,-77.5,-214,-77.5</points>
<connection>
<GID>359</GID>
<name>IN_B_1</name></connection>
<intersection>-239 10</intersection>
<intersection>-233 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-233,-77.5,-233,-62.5</points>
<intersection>-77.5 1</intersection>
<intersection>-62.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-233,-62.5,-190,-62.5</points>
<connection>
<GID>358</GID>
<name>IN_B_1</name></connection>
<intersection>-233 8</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-239,-82,-239,-77.5</points>
<intersection>-82 14</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-241,-82,-239,-82</points>
<connection>
<GID>345</GID>
<name>OUT_1</name></connection>
<intersection>-239 10</intersection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-235.5,-79.5,-214,-79.5</points>
<connection>
<GID>359</GID>
<name>IN_B_3</name></connection>
<intersection>-235.5 8</intersection>
<intersection>-230.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-230.5,-79.5,-230.5,-64.5</points>
<intersection>-79.5 1</intersection>
<intersection>-64.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-230.5,-64.5,-190,-64.5</points>
<connection>
<GID>358</GID>
<name>IN_B_3</name></connection>
<intersection>-230.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-235.5,-84,-235.5,-79.5</points>
<intersection>-84 9</intersection>
<intersection>-79.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-241,-84,-235.5,-84</points>
<connection>
<GID>345</GID>
<name>OUT_3</name></connection>
<intersection>-235.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-214.5,-86.5,-214,-86.5</points>
<connection>
<GID>361</GID>
<name>OUT_0</name></connection>
<connection>
<GID>359</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249.5,-50.5,-249.5,-46.5</points>
<intersection>-50.5 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-298.5,-50.5,-249.5,-50.5</points>
<intersection>-298.5 3</intersection>
<intersection>-249.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-249.5,-46.5,-249,-46.5</points>
<connection>
<GID>343</GID>
<name>IN_2</name></connection>
<intersection>-249.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-298.5,-53,-298.5,-50.5</points>
<connection>
<GID>339</GID>
<name>OUT_2</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-298.5,-53,-249,-53</points>
<intersection>-298.5 3</intersection>
<intersection>-249 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-249,-53,-249,-47.5</points>
<connection>
<GID>343</GID>
<name>IN_3</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>-298.5,-53,-298.5,-51</points>
<connection>
<GID>339</GID>
<name>OUT_3</name></connection>
<intersection>-53 1</intersection></vsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-162.5,-79,-162.5,-79</points>
<connection>
<GID>362</GID>
<name>N_in2</name></connection>
<connection>
<GID>369</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-162.5,-81,-162.5,-81</points>
<connection>
<GID>369</GID>
<name>N_in2</name></connection>
<connection>
<GID>370</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-246,-67,-246,-50.5</points>
<connection>
<GID>343</GID>
<name>carry_out</name></connection>
<connection>
<GID>386</GID>
<name>IN_1</name></connection>
<intersection>-57 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-246,-57,-237,-57</points>
<connection>
<GID>377</GID>
<name>IN_1</name></connection>
<intersection>-246 0</intersection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-167,-31,-167,-28</points>
<connection>
<GID>363</GID>
<name>IN_3</name></connection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-31,-167,-31</points>
<connection>
<GID>346</GID>
<name>OUT_3</name></connection>
<intersection>-167 0</intersection></hsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-167,-30,-167,-29</points>
<connection>
<GID>363</GID>
<name>IN_2</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-30,-167,-30</points>
<connection>
<GID>346</GID>
<name>OUT_2</name></connection>
<intersection>-167 0</intersection></hsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-167,-30,-167,-29</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<intersection>-29 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-182,-29,-167,-29</points>
<connection>
<GID>346</GID>
<name>OUT_1</name></connection>
<intersection>-167 3</intersection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-167,-31,-167,-28</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-28,-167,-28</points>
<connection>
<GID>346</GID>
<name>OUT_0</name></connection>
<intersection>-167 0</intersection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-210,-54.5,-207.5,-54.5</points>
<intersection>-210 6</intersection>
<intersection>-207.5 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-210,-54.5,-210,-54</points>
<connection>
<GID>350</GID>
<name>A_less_B</name></connection>
<intersection>-54.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-207.5,-54.5,-207.5,-54</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-54.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-165.5,-68,-165.5,-65</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-65,-165.5,-65</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>-165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-182.5,-67,-182.5,-66</points>
<intersection>-67 1</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182.5,-67,-165.5,-67</points>
<connection>
<GID>365</GID>
<name>IN_1</name></connection>
<intersection>-182.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-182.5,-66,-182,-66</points>
<connection>
<GID>358</GID>
<name>OUT_1</name></connection>
<intersection>-182.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-165.5,-67,-165.5,-66</points>
<connection>
<GID>365</GID>
<name>IN_2</name></connection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-67,-165.5,-67</points>
<connection>
<GID>358</GID>
<name>OUT_2</name></connection>
<intersection>-165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-165,-68,-165,-65</points>
<intersection>-68 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-68,-165,-68</points>
<connection>
<GID>358</GID>
<name>OUT_3</name></connection>
<intersection>-165 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-165.5,-65,-165,-65</points>
<connection>
<GID>365</GID>
<name>IN_3</name></connection>
<intersection>-165 0</intersection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>533,-16,533,-15</points>
<connection>
<GID>311</GID>
<name>load</name></connection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>533.5,-15,533.5,-14.5</points>
<connection>
<GID>413</GID>
<name>OUT_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>533,-15,533.5,-15</points>
<intersection>533 0</intersection>
<intersection>533.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-163,-83,-162.5,-83</points>
<connection>
<GID>371</GID>
<name>N_in3</name></connection>
<connection>
<GID>370</GID>
<name>N_in2</name></connection>
<intersection>-163 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-163,-83,-163,-82</points>
<intersection>-83 1</intersection>
<intersection>-82 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-163.5,-82,-163,-82</points>
<connection>
<GID>370</GID>
<name>N_in0</name></connection>
<intersection>-163 4</intersection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-187,-58.5,-187,-37.5</points>
<connection>
<GID>346</GID>
<name>carry_out</name></connection>
<connection>
<GID>358</GID>
<name>carry_in</name></connection>
<intersection>-58.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-225,-58.5,-187,-58.5</points>
<intersection>-225 9</intersection>
<intersection>-187 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-225,-84.5,-225,-58.5</points>
<intersection>-84.5 10</intersection>
<intersection>-58.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-225,-84.5,-220,-84.5</points>
<connection>
<GID>367</GID>
<name>IN_1</name></connection>
<intersection>-225 9</intersection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-220,-82.5,-220,-82.5</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>567,-33.5,567,2</points>
<intersection>-33.5 5</intersection>
<intersection>2 13</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>524.5,-33.5,584,-33.5</points>
<connection>
<GID>310</GID>
<name>IN_7</name></connection>
<intersection>524.5 8</intersection>
<intersection>567 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>524.5,-33.5,524.5,-17</points>
<intersection>-33.5 5</intersection>
<intersection>-17 14</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>553.5,2,567,2</points>
<connection>
<GID>412</GID>
<name>OUT_3</name></connection>
<intersection>567 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>524.5,-17,530,-17</points>
<intersection>524.5 8</intersection>
<intersection>530 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>530,-18,530,-17</points>
<connection>
<GID>311</GID>
<name>IN_7</name></connection>
<intersection>-17 14</intersection></vsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-157,-77,-157,-13</points>
<intersection>-77 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-244,-13,-157,-13</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<intersection>-157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-162.5,-77,-157,-77</points>
<connection>
<GID>362</GID>
<name>N_in3</name></connection>
<intersection>-157 0</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-206.5,-48,-206.5,-35.5</points>
<connection>
<GID>364</GID>
<name>OUT</name></connection>
<intersection>-39.5 21</intersection>
<intersection>-35.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-206.5,-35.5,-197.5,-35.5</points>
<connection>
<GID>374</GID>
<name>IN_1</name></connection>
<intersection>-206.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-206.5,-39.5,-197.5,-39.5</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<intersection>-206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-190.5,-38.5,-190.5,-33.5</points>
<intersection>-38.5 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-190.5,-33.5,-190,-33.5</points>
<connection>
<GID>346</GID>
<name>IN_2</name></connection>
<intersection>-190.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-191.5,-38.5,-190.5,-38.5</points>
<connection>
<GID>375</GID>
<name>OUT</name></connection>
<intersection>-190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-191,-34.5,-191,-32.5</points>
<intersection>-34.5 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-191,-32.5,-190,-32.5</points>
<connection>
<GID>346</GID>
<name>IN_1</name></connection>
<intersection>-191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-191.5,-34.5,-191,-34.5</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<intersection>-191 0</intersection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-191,-31.5,-191,-30.5</points>
<intersection>-31.5 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-191,-31.5,-190,-31.5</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>-191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-191.5,-30.5,-191,-30.5</points>
<connection>
<GID>373</GID>
<name>OUT</name></connection>
<intersection>-191 0</intersection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-190,-42.5,-190,-34.5</points>
<connection>
<GID>346</GID>
<name>IN_3</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-191.5,-42.5,-190,-42.5</points>
<connection>
<GID>376</GID>
<name>OUT</name></connection>
<intersection>-190 0</intersection></hsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-197.5,-31.5,-197.5,-31.5</points>
<connection>
<GID>373</GID>
<name>IN_1</name></connection>
<connection>
<GID>379</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-197.5,-43.5,-197.5,-43.5</points>
<connection>
<GID>376</GID>
<name>IN_1</name></connection>
<connection>
<GID>380</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-199.5,-89.5,-199.5,-71.5</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>-75.5 21</intersection>
<intersection>-71.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-199.5,-71.5,-197,-71.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>-199.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-199.5,-75.5,-197,-75.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>-199.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-197,-67.5,-197,-67.5</points>
<connection>
<GID>336</GID>
<name>IN_1</name></connection>
<connection>
<GID>381</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-197,-79.5,-197,-79.5</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<connection>
<GID>341</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-270.5,-79.5,-270.5,-18.5</points>
<intersection>-79.5 246</intersection>
<intersection>-75.5 247</intersection>
<intersection>-71.5 248</intersection>
<intersection>-67.5 249</intersection>
<intersection>-38.5 101</intersection>
<intersection>-34.5 39</intersection>
<intersection>-30.5 29</intersection>
<intersection>-26.5 28</intersection>
<intersection>-18.5 30</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-270.5,-26.5,-266,-26.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-270.5,-30.5,-266,-30.5</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-270.5,-18.5,-187,-18.5</points>
<connection>
<GID>356</GID>
<name>OUT</name></connection>
<intersection>-270.5 0</intersection>
<intersection>-244 233</intersection>
<intersection>-202 37</intersection>
<intersection>-187 226</intersection></hsegment>
<vsegment>
<ID>37</ID>
<points>-202,-95.5,-202,-18.5</points>
<intersection>-95.5 255</intersection>
<intersection>-77.5 90</intersection>
<intersection>-73.5 98</intersection>
<intersection>-69.5 95</intersection>
<intersection>-65.5 96</intersection>
<intersection>-41.5 237</intersection>
<intersection>-37.5 48</intersection>
<intersection>-33.5 45</intersection>
<intersection>-29.5 228</intersection>
<intersection>-18.5 30</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>-270.5,-34.5,-266,-34.5</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>-202,-33.5,-197.5,-33.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-202,-37.5,-197.5,-37.5</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>90</ID>
<points>-202,-77.5,-197,-77.5</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>95</ID>
<points>-202,-69.5,-197,-69.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>96</ID>
<points>-202,-65.5,-197,-65.5</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>98</ID>
<points>-202,-73.5,-197,-73.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>101</ID>
<points>-270.5,-38.5,-266,-38.5</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<vsegment>
<ID>226</ID>
<points>-187,-21.5,-187,-18.5</points>
<connection>
<GID>346</GID>
<name>carry_in</name></connection>
<intersection>-18.5 30</intersection></vsegment>
<hsegment>
<ID>228</ID>
<points>-202,-29.5,-197.5,-29.5</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<vsegment>
<ID>233</ID>
<points>-244,-67,-244,-18.5</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>-55 234</intersection>
<intersection>-34.5 256</intersection>
<intersection>-18.5 30</intersection></vsegment>
<hsegment>
<ID>234</ID>
<points>-244,-55,-237,-55</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>-244 233</intersection></hsegment>
<hsegment>
<ID>237</ID>
<points>-202,-41.5,-197.5,-41.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>246</ID>
<points>-270.5,-79.5,-267,-79.5</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>247</ID>
<points>-270.5,-75.5,-267,-75.5</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>248</ID>
<points>-270.5,-71.5,-267,-71.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>249</ID>
<points>-270.5,-67.5,-267,-67.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>255</ID>
<points>-202,-95.5,-200.5,-95.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>256</ID>
<points>-246,-34.5,-244,-34.5</points>
<connection>
<GID>343</GID>
<name>carry_in</name></connection>
<intersection>-244 233</intersection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-190,-78.5,-190,-71.5</points>
<connection>
<GID>358</GID>
<name>IN_3</name></connection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-191,-78.5,-190,-78.5</points>
<connection>
<GID>341</GID>
<name>OUT</name></connection>
<intersection>-190 0</intersection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-190.5,-68.5,-190.5,-66.5</points>
<intersection>-68.5 1</intersection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-190.5,-68.5,-190,-68.5</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>-190.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-191,-66.5,-190.5,-66.5</points>
<connection>
<GID>336</GID>
<name>OUT</name></connection>
<intersection>-190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-191,-70.5,-191,-69.5</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-191,-69.5,-190,-69.5</points>
<connection>
<GID>358</GID>
<name>IN_1</name></connection>
<intersection>-191 0</intersection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-190.5,-74.5,-190.5,-70.5</points>
<intersection>-74.5 4</intersection>
<intersection>-70.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-190.5,-70.5,-190,-70.5</points>
<connection>
<GID>358</GID>
<name>IN_2</name></connection>
<intersection>-190.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-191,-74.5,-190.5,-74.5</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<intersection>-190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,-40.5,-268,-34</points>
<intersection>-40.5 5</intersection>
<intersection>-34 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-272,-34,-268,-34</points>
<connection>
<GID>335</GID>
<name>OUT_3</name></connection>
<intersection>-268 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-268,-40.5,-266,-40.5</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,-36.5,-268,-36</points>
<intersection>-36.5 5</intersection>
<intersection>-36 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-272,-36,-268,-36</points>
<connection>
<GID>335</GID>
<name>OUT_2</name></connection>
<intersection>-268 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-268,-36.5,-266,-36.5</points>
<connection>
<GID>357</GID>
<name>IN_1</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,-38,-268,-32.5</points>
<intersection>-38 4</intersection>
<intersection>-32.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-272,-38,-268,-38</points>
<connection>
<GID>335</GID>
<name>OUT_1</name></connection>
<intersection>-268 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-268,-32.5,-266,-32.5</points>
<connection>
<GID>348</GID>
<name>IN_1</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,-40,-268,-28.5</points>
<intersection>-40 4</intersection>
<intersection>-28.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-272,-40,-268,-40</points>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection>
<intersection>-268 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-268,-28.5,-266,-28.5</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-269,-81.5,-269,-75</points>
<intersection>-81.5 3</intersection>
<intersection>-75 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-269,-81.5,-267,-81.5</points>
<connection>
<GID>334</GID>
<name>IN_1</name></connection>
<intersection>-269 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-273.5,-75,-269,-75</points>
<connection>
<GID>342</GID>
<name>OUT_3</name></connection>
<intersection>-269 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-269,-77.5,-269,-77</points>
<intersection>-77.5 3</intersection>
<intersection>-77 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-269,-77.5,-267,-77.5</points>
<connection>
<GID>333</GID>
<name>IN_1</name></connection>
<intersection>-269 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-273.5,-77,-269,-77</points>
<connection>
<GID>342</GID>
<name>OUT_2</name></connection>
<intersection>-269 0</intersection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-269,-79,-269,-73.5</points>
<intersection>-79 4</intersection>
<intersection>-73.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-269,-73.5,-267,-73.5</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<intersection>-269 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-273.5,-79,-269,-79</points>
<connection>
<GID>342</GID>
<name>OUT_1</name></connection>
<intersection>-269 0</intersection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-269,-81,-269,-69.5</points>
<intersection>-81 4</intersection>
<intersection>-69.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-269,-69.5,-267,-69.5</points>
<connection>
<GID>331</GID>
<name>IN_1</name></connection>
<intersection>-269 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-273.5,-81,-269,-81</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<intersection>-269 0</intersection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-246,-98.5,-246,-90.5</points>
<connection>
<GID>345</GID>
<name>carry_out</name></connection>
<intersection>-98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-246,-98.5,-206.5,-98.5</points>
<connection>
<GID>366</GID>
<name>IN_1</name></connection>
<intersection>-246 0</intersection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-254.5,-37.5,-254.5,-27.5</points>
<intersection>-37.5 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-254.5,-37.5,-249,-37.5</points>
<connection>
<GID>343</GID>
<name>IN_B_0</name></connection>
<intersection>-254.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-260,-27.5,-254.5,-27.5</points>
<connection>
<GID>347</GID>
<name>OUT</name></connection>
<intersection>-254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-254.5,-38.5,-254.5,-31.5</points>
<intersection>-38.5 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-260,-31.5,-254.5,-31.5</points>
<connection>
<GID>348</GID>
<name>OUT</name></connection>
<intersection>-254.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-254.5,-38.5,-249,-38.5</points>
<connection>
<GID>343</GID>
<name>IN_B_1</name></connection>
<intersection>-254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-254.5,-39.5,-254.5,-35.5</points>
<intersection>-39.5 1</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-254.5,-39.5,-249,-39.5</points>
<connection>
<GID>343</GID>
<name>IN_B_2</name></connection>
<intersection>-254.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-260,-35.5,-254.5,-35.5</points>
<connection>
<GID>357</GID>
<name>OUT</name></connection>
<intersection>-254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-254.5,-40.5,-254.5,-39.5</points>
<intersection>-40.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-260,-39.5,-254.5,-39.5</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<intersection>-254.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-254.5,-40.5,-249,-40.5</points>
<connection>
<GID>343</GID>
<name>IN_B_3</name></connection>
<intersection>-254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-255,-77.5,-255,-68.5</points>
<intersection>-77.5 1</intersection>
<intersection>-68.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-255,-77.5,-249,-77.5</points>
<connection>
<GID>345</GID>
<name>IN_B_0</name></connection>
<intersection>-255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-261,-68.5,-255,-68.5</points>
<connection>
<GID>331</GID>
<name>OUT</name></connection>
<intersection>-255 0</intersection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-255,-78.5,-255,-72.5</points>
<intersection>-78.5 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-261,-72.5,-255,-72.5</points>
<connection>
<GID>332</GID>
<name>OUT</name></connection>
<intersection>-255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-255,-78.5,-249,-78.5</points>
<connection>
<GID>345</GID>
<name>IN_B_1</name></connection>
<intersection>-255 0</intersection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-255,-79.5,-255,-76.5</points>
<intersection>-79.5 1</intersection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-255,-79.5,-249,-79.5</points>
<connection>
<GID>345</GID>
<name>IN_B_2</name></connection>
<intersection>-255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-261,-76.5,-255,-76.5</points>
<connection>
<GID>333</GID>
<name>OUT</name></connection>
<intersection>-255 0</intersection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-261,-80.5,-249,-80.5</points>
<connection>
<GID>334</GID>
<name>OUT</name></connection>
<connection>
<GID>345</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-205.5,-56,-205.5,-54</points>
<connection>
<GID>364</GID>
<name>IN_1</name></connection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-231,-56,-205.5,-56</points>
<connection>
<GID>377</GID>
<name>OUT</name></connection>
<intersection>-205.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>564.5,-34.5,564.5,3</points>
<intersection>-34.5 1</intersection>
<intersection>3 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-34.5,584,-34.5</points>
<connection>
<GID>310</GID>
<name>IN_6</name></connection>
<intersection>527.5 6</intersection>
<intersection>564.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>527.5,-34.5,527.5,-19</points>
<intersection>-34.5 1</intersection>
<intersection>-19 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>553.5,3,564.5,3</points>
<connection>
<GID>412</GID>
<name>OUT_2</name></connection>
<intersection>564.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>527.5,-19,530,-19</points>
<connection>
<GID>311</GID>
<name>IN_6</name></connection>
<intersection>527.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-214,-83.5,-214,-83.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-198.5,-97.5,-198.5,-95.5</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-200.5,-97.5,-198.5,-97.5</points>
<connection>
<GID>366</GID>
<name>OUT</name></connection>
<intersection>-198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>561.5,-35.5,561.5,4</points>
<intersection>-35.5 1</intersection>
<intersection>4 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>526.5,-35.5,584,-35.5</points>
<connection>
<GID>310</GID>
<name>IN_5</name></connection>
<intersection>526.5 6</intersection>
<intersection>561.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>526.5,-35.5,526.5,-20</points>
<intersection>-35.5 1</intersection>
<intersection>-20 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>553.5,4,561.5,4</points>
<connection>
<GID>412</GID>
<name>OUT_1</name></connection>
<intersection>561.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>526.5,-20,530,-20</points>
<connection>
<GID>311</GID>
<name>IN_5</name></connection>
<intersection>526.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-172,-78,-172,-77.5</points>
<connection>
<GID>385</GID>
<name>N_in3</name></connection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-187,-78,-172,-78</points>
<intersection>-187 2</intersection>
<intersection>-172 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-187,-78,-187,-74.5</points>
<connection>
<GID>358</GID>
<name>carry_out</name></connection>
<intersection>-78 1</intersection></vsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>558.5,-36.5,558.5,5</points>
<intersection>-36.5 1</intersection>
<intersection>5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>529,-36.5,584,-36.5</points>
<connection>
<GID>310</GID>
<name>IN_4</name></connection>
<intersection>529 6</intersection>
<intersection>558.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>529,-36.5,529,-21</points>
<intersection>-36.5 1</intersection>
<intersection>-21 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>553.5,5,558.5,5</points>
<connection>
<GID>412</GID>
<name>OUT_0</name></connection>
<intersection>558.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>529,-21,530,-21</points>
<connection>
<GID>311</GID>
<name>IN_4</name></connection>
<intersection>529 6</intersection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>572.5,-37.5,572.5,24</points>
<intersection>-37.5 1</intersection>
<intersection>24 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>529.5,-37.5,584,-37.5</points>
<connection>
<GID>310</GID>
<name>IN_3</name></connection>
<intersection>529.5 6</intersection>
<intersection>572.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>529.5,-37.5,529.5,-22</points>
<intersection>-37.5 1</intersection>
<intersection>-22 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>553.5,24,572.5,24</points>
<connection>
<GID>411</GID>
<name>OUT_3</name></connection>
<intersection>572.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>529.5,-22,530,-22</points>
<connection>
<GID>311</GID>
<name>IN_3</name></connection>
<intersection>529.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-208,-96.5,-208,-89.5</points>
<connection>
<GID>359</GID>
<name>A_less_B</name></connection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-208,-96.5,-206.5,-96.5</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>-208 0</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-162.5,-84,-162.5,-80</points>
<intersection>-84 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-162.5,-84,-161.5,-84</points>
<connection>
<GID>371</GID>
<name>N_in1</name></connection>
<intersection>-162.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-163.5,-80,-162.5,-80</points>
<connection>
<GID>369</GID>
<name>N_in0</name></connection>
<intersection>-162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-245,-74.5,-245,-73</points>
<connection>
<GID>386</GID>
<name>OUT</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-246,-74.5,-245,-74.5</points>
<connection>
<GID>345</GID>
<name>carry_in</name></connection>
<intersection>-245 0</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-81.5,359,-78</points>
<connection>
<GID>302</GID>
<name>OUT_3</name></connection>
<intersection>-81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-81.5,364,-81.5</points>
<connection>
<GID>308</GID>
<name>IN_3</name></connection>
<intersection>359 0</intersection></hsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>360,-82.5,360,-78</points>
<connection>
<GID>302</GID>
<name>OUT_2</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360,-82.5,364,-82.5</points>
<connection>
<GID>308</GID>
<name>IN_2</name></connection>
<intersection>360 0</intersection></hsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361,-83.5,361,-78</points>
<connection>
<GID>302</GID>
<name>OUT_1</name></connection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361,-83.5,364,-83.5</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>361 0</intersection></hsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362,-84.5,362,-78</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>362,-84.5,364,-84.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>362 0</intersection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>314.5,-58.5,339,-58.5</points>
<intersection>314.5 26</intersection>
<intersection>327 39</intersection>
<intersection>331 27</intersection>
<intersection>335 28</intersection>
<intersection>339 29</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>314.5,-82.5,314.5,-56.5</points>
<connection>
<GID>397</GID>
<name>OUT_0</name></connection>
<intersection>-82.5 40</intersection>
<intersection>-69 30</intersection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>331,-60,331,-58.5</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>335,-60,335,-58.5</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>339,-60,339,-58.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>314.5,-69,324,-69</points>
<intersection>314.5 26</intersection>
<intersection>322 42</intersection>
<intersection>324 32</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>324,-70,324,-69</points>
<connection>
<GID>391</GID>
<name>IN_1</name></connection>
<intersection>-69 30</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>327,-60,327,-58.5</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>40</ID>
<points>314.5,-82.5,317,-82.5</points>
<connection>
<GID>396</GID>
<name>N_in0</name></connection>
<intersection>314.5 26</intersection></hsegment>
<vsegment>
<ID>42</ID>
<points>322,-70,322,-69</points>
<connection>
<GID>391</GID>
<name>IN_3</name></connection>
<intersection>-69 30</intersection></vsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334.5,-69,334.5,-66.5</points>
<intersection>-69 3</intersection>
<intersection>-66.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>338,-66.5,338,-66</points>
<connection>
<GID>390</GID>
<name>OUT</name></connection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>334.5,-66.5,338,-66.5</points>
<intersection>334.5 0</intersection>
<intersection>338 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>332,-69,334.5,-69</points>
<intersection>332 4</intersection>
<intersection>334.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>332,-70,332,-69</points>
<connection>
<GID>391</GID>
<name>IN_B_0</name></connection>
<intersection>-69 3</intersection></vsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331,-70,331,-68.5</points>
<connection>
<GID>391</GID>
<name>IN_B_1</name></connection>
<intersection>-68.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>334,-68.5,334,-66</points>
<connection>
<GID>389</GID>
<name>OUT</name></connection>
<intersection>-68.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>331,-68.5,334,-68.5</points>
<intersection>331 0</intersection>
<intersection>334 1</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,-70,330,-66</points>
<connection>
<GID>388</GID>
<name>OUT</name></connection>
<connection>
<GID>391</GID>
<name>IN_B_2</name></connection></vsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327.5,-69,327.5,-66</points>
<intersection>-69 3</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>326,-66,327.5,-66</points>
<connection>
<GID>387</GID>
<name>OUT</name></connection>
<intersection>327.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>327.5,-69,329,-69</points>
<intersection>327.5 0</intersection>
<intersection>329 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>329,-70,329,-69</points>
<connection>
<GID>391</GID>
<name>IN_B_3</name></connection>
<intersection>-69 3</intersection></vsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323,-82.5,323,-82.5</points>
<connection>
<GID>393</GID>
<name>N_in0</name></connection>
<connection>
<GID>394</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321,-82.5,321,-82.5</points>
<connection>
<GID>394</GID>
<name>N_in0</name></connection>
<connection>
<GID>395</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319,-82.5,319,-82.5</points>
<connection>
<GID>395</GID>
<name>N_in0</name></connection>
<connection>
<GID>396</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325.5,-81.5,325.5,-78</points>
<connection>
<GID>391</GID>
<name>OUT_3</name></connection>
<intersection>-81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>325.5,-81.5,330.5,-81.5</points>
<connection>
<GID>392</GID>
<name>IN_3</name></connection>
<intersection>325.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326.5,-82.5,326.5,-78</points>
<connection>
<GID>391</GID>
<name>OUT_2</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>326.5,-82.5,330.5,-82.5</points>
<connection>
<GID>392</GID>
<name>IN_2</name></connection>
<intersection>326.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327.5,-83.5,327.5,-78</points>
<connection>
<GID>391</GID>
<name>OUT_1</name></connection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>327.5,-83.5,330.5,-83.5</points>
<connection>
<GID>392</GID>
<name>IN_1</name></connection>
<intersection>327.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328.5,-84.5,328.5,-78</points>
<connection>
<GID>391</GID>
<name>OUT_0</name></connection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>328.5,-84.5,330.5,-84.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>328.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-60,337,-57</points>
<connection>
<GID>390</GID>
<name>IN_1</name></connection>
<connection>
<GID>297</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,-60,333,-58</points>
<connection>
<GID>389</GID>
<name>IN_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>336,-58,336,-57</points>
<connection>
<GID>297</GID>
<name>OUT_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>333,-58,336,-58</points>
<intersection>333 0</intersection>
<intersection>336 1</intersection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329,-60,329,-58</points>
<connection>
<GID>388</GID>
<name>IN_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>335,-58,335,-57</points>
<connection>
<GID>297</GID>
<name>OUT_2</name></connection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>329,-58,335,-58</points>
<intersection>329 0</intersection>
<intersection>335 1</intersection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,-57.5,334,-57</points>
<connection>
<GID>297</GID>
<name>OUT_3</name></connection>
<intersection>-57.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>325,-60,325,-57.5</points>
<connection>
<GID>387</GID>
<name>IN_1</name></connection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>325,-57.5,334,-57.5</points>
<intersection>325 1</intersection>
<intersection>334 0</intersection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326,-40,326,-40</points>
<connection>
<GID>398</GID>
<name>OUT</name></connection>
<connection>
<GID>290</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325,-34,325,-34</points>
<connection>
<GID>398</GID>
<name>IN_1</name></connection>
<connection>
<GID>399</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>574,-38.5,574,25</points>
<intersection>-38.5 1</intersection>
<intersection>25 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>530,-38.5,584,-38.5</points>
<connection>
<GID>310</GID>
<name>IN_2</name></connection>
<intersection>530 6</intersection>
<intersection>574 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>530,-38.5,530,-23</points>
<connection>
<GID>311</GID>
<name>IN_2</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>553.5,25,574,25</points>
<connection>
<GID>411</GID>
<name>OUT_2</name></connection>
<intersection>574 0</intersection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350,-46.5,351.5,-46.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<connection>
<GID>284</GID>
<name>A_less_B</name></connection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>343.5,-52,359,-52</points>
<connection>
<GID>288</GID>
<name>carry_out</name></connection>
<intersection>343.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>343.5,-52,343.5,-38.5</points>
<connection>
<GID>297</GID>
<name>carry_in</name></connection>
<intersection>-52 1</intersection>
<intersection>-38.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>329,-38.5,343.5,-38.5</points>
<intersection>329 5</intersection>
<intersection>343.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>329,-38.5,329,-34</points>
<intersection>-38.5 4</intersection>
<intersection>-34 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>327,-34,329,-34</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>329 5</intersection></hsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>575.5,-39.5,575.5,26</points>
<intersection>-39.5 1</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>528,-39.5,584,-39.5</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<intersection>528 8</intersection>
<intersection>575.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>553.5,26,575.5,26</points>
<connection>
<GID>411</GID>
<name>OUT_1</name></connection>
<intersection>575.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>528,-39.5,528,-24</points>
<intersection>-39.5 1</intersection>
<intersection>-24 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>528,-24,530,-24</points>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<intersection>528 8</intersection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>577,-40.5,577,27</points>
<intersection>-40.5 1</intersection>
<intersection>27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525.5,-40.5,584,-40.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>525.5 7</intersection>
<intersection>577 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>553.5,27,577,27</points>
<connection>
<GID>411</GID>
<name>OUT_0</name></connection>
<intersection>577 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>525.5,-40.5,525.5,-25</points>
<intersection>-40.5 1</intersection>
<intersection>-25 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>525.5,-25,530,-25</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>525.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>548.5,11.5,548.5,17.5</points>
<connection>
<GID>412</GID>
<name>carry_in</name></connection>
<connection>
<GID>411</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515,-32.5,515,5</points>
<connection>
<GID>673</GID>
<name>OUT_0</name></connection>
<intersection>-28.5 16</intersection>
<intersection>-12 6</intersection>
<intersection>5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>510,5,516,5</points>
<connection>
<GID>313</GID>
<name>clear</name></connection>
<intersection>515 0</intersection>
<intersection>516 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>510,-12,515,-12</points>
<intersection>510 13</intersection>
<intersection>515 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>516,5,516,22</points>
<intersection>5 5</intersection>
<intersection>22 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>511,22,516,22</points>
<connection>
<GID>312</GID>
<name>clear</name></connection>
<intersection>516 7</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>510,-12,510,-11</points>
<connection>
<GID>325</GID>
<name>clear</name></connection>
<intersection>-12 6</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>515,-28.5,535,-28.5</points>
<intersection>515 0</intersection>
<intersection>535 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>535,-28.5,535,-27</points>
<connection>
<GID>311</GID>
<name>clear</name></connection>
<intersection>-28.5 16</intersection></vsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>501,24.5,501,28.5</points>
<intersection>24.5 2</intersection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>501,28.5,507.5,28.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>501 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>495,24.5,501,24.5</points>
<connection>
<GID>223</GID>
<name>OUT_3</name></connection>
<intersection>501 0</intersection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502,22.5,502,27.5</points>
<intersection>22.5 2</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>502,27.5,507.5,27.5</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<intersection>502 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>495,22.5,502,22.5</points>
<connection>
<GID>223</GID>
<name>OUT_2</name></connection>
<intersection>502 0</intersection></hsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502,20.5,502,26.5</points>
<intersection>20.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>495,20.5,502,20.5</points>
<connection>
<GID>223</GID>
<name>OUT_1</name></connection>
<intersection>502 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>502,26.5,507.5,26.5</points>
<connection>
<GID>312</GID>
<name>IN_2</name></connection>
<intersection>502 0</intersection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>503.5,18.5,503.5,25.5</points>
<intersection>18.5 1</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>495,18.5,503.5,18.5</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>503.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503.5,25.5,507.5,25.5</points>
<connection>
<GID>312</GID>
<name>IN_3</name></connection>
<intersection>503.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>501,8,501,8.5</points>
<intersection>8 2</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>501,8.5,506.5,8.5</points>
<connection>
<GID>313</GID>
<name>IN_3</name></connection>
<intersection>501 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>494.5,8,501,8</points>
<connection>
<GID>260</GID>
<name>OUT_3</name></connection>
<intersection>501 0</intersection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502,6,502,9.5</points>
<intersection>6 2</intersection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>502,9.5,506.5,9.5</points>
<connection>
<GID>313</GID>
<name>IN_2</name></connection>
<intersection>502 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>494.5,6,502,6</points>
<connection>
<GID>260</GID>
<name>OUT_2</name></connection>
<intersection>502 0</intersection></hsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>503,4,503,10.5</points>
<intersection>4 2</intersection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503,10.5,506.5,10.5</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>503 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>494.5,4,503,4</points>
<connection>
<GID>260</GID>
<name>OUT_1</name></connection>
<intersection>503 0</intersection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>498.5,2,498.5,14</points>
<intersection>2 2</intersection>
<intersection>14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>498.5,14,506.5,14</points>
<intersection>498.5 0</intersection>
<intersection>506.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>494.5,2,498.5,2</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<intersection>498.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>506.5,11.5,506.5,14</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>14 1</intersection></vsegment></shape></wire>
<wire>
<ID>768</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,15,510,15.5</points>
<connection>
<GID>313</GID>
<name>shift_enable</name></connection>
<intersection>15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>509.5,15.5,509.5,16</points>
<connection>
<GID>383</GID>
<name>OUT_0</name></connection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>509.5,15.5,510,15.5</points>
<intersection>509.5 1</intersection>
<intersection>510 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-22.5313,2284.15,1755.47,1357.15</PageViewport></page 3>
<page 4>
<PageViewport>365.559,1998.87,543.56,1906.07</PageViewport>
<gate>
<ID>585</ID>
<type>DD_KEYPAD_HEX</type>
<position>491.5,1937</position>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>414</ID>
<type>DA_FROM</type>
<position>406.5,1963</position>
<input>
<ID>IN_0</ID>603 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>417</ID>
<type>DA_FROM</type>
<position>406.5,1965</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>422</ID>
<type>DA_FROM</type>
<position>406.5,1967</position>
<input>
<ID>IN_0</ID>604 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>424</ID>
<type>DA_FROM</type>
<position>406.5,1969</position>
<input>
<ID>IN_0</ID>622 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>425</ID>
<type>DA_FROM</type>
<position>406.5,1971</position>
<input>
<ID>IN_0</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>427</ID>
<type>DA_FROM</type>
<position>406.5,1973</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>430</ID>
<type>DA_FROM</type>
<position>406.5,1975</position>
<input>
<ID>IN_0</ID>606 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>431</ID>
<type>DA_FROM</type>
<position>406.5,1977</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>432</ID>
<type>DA_FROM</type>
<position>406.5,1979</position>
<input>
<ID>IN_0</ID>612 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>433</ID>
<type>AE_REGISTER8</type>
<position>441,1962.5</position>
<input>
<ID>IN_0</ID>628 </input>
<input>
<ID>IN_1</ID>627 </input>
<input>
<ID>IN_2</ID>626 </input>
<input>
<ID>IN_3</ID>625 </input>
<output>
<ID>OUT_0</ID>716 </output>
<output>
<ID>OUT_1</ID>717 </output>
<output>
<ID>OUT_2</ID>718 </output>
<output>
<ID>OUT_3</ID>719 </output>
<input>
<ID>clock</ID>738 </input>
<input>
<ID>load</ID>738 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>434</ID>
<type>AE_OR2</type>
<position>461,1934</position>
<input>
<ID>IN_0</ID>746 </input>
<input>
<ID>IN_1</ID>745 </input>
<output>
<ID>OUT</ID>744 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>435</ID>
<type>DA_FROM</type>
<position>460,1929</position>
<input>
<ID>IN_0</ID>746 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>436</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>433,1970</position>
<input>
<ID>IN_0</ID>615 </input>
<input>
<ID>IN_1</ID>616 </input>
<input>
<ID>IN_2</ID>620 </input>
<input>
<ID>IN_3</ID>619 </input>
<output>
<ID>OUT_0</ID>628 </output>
<output>
<ID>OUT_1</ID>627 </output>
<output>
<ID>OUT_2</ID>626 </output>
<output>
<ID>OUT_3</ID>625 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>437</ID>
<type>DE_OR8</type>
<position>422,1959</position>
<input>
<ID>IN_0</ID>614 </input>
<input>
<ID>IN_1</ID>614 </input>
<input>
<ID>IN_2</ID>614 </input>
<input>
<ID>IN_3</ID>612 </input>
<input>
<ID>IN_4</ID>603 </input>
<input>
<ID>IN_5</ID>604 </input>
<input>
<ID>IN_6</ID>605 </input>
<input>
<ID>IN_7</ID>606 </input>
<output>
<ID>OUT</ID>615 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>438</ID>
<type>FF_GND</type>
<position>418,1960.5</position>
<output>
<ID>OUT_0</ID>614 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>439</ID>
<type>AE_OR2</type>
<position>422,1981</position>
<input>
<ID>IN_0</ID>612 </input>
<input>
<ID>IN_1</ID>621 </input>
<output>
<ID>OUT</ID>619 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>440</ID>
<type>AE_OR4</type>
<position>421,1967</position>
<input>
<ID>IN_0</ID>606 </input>
<input>
<ID>IN_1</ID>618 </input>
<input>
<ID>IN_2</ID>604 </input>
<input>
<ID>IN_3</ID>617 </input>
<output>
<ID>OUT</ID>616 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>441</ID>
<type>AE_OR4</type>
<position>421,1975</position>
<input>
<ID>IN_0</ID>606 </input>
<input>
<ID>IN_1</ID>618 </input>
<input>
<ID>IN_2</ID>605 </input>
<input>
<ID>IN_3</ID>622 </input>
<output>
<ID>OUT</ID>620 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>444</ID>
<type>DA_FROM</type>
<position>406.5,1961</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>471</ID>
<type>AE_OR4</type>
<position>430,1959</position>
<input>
<ID>IN_0</ID>619 </input>
<input>
<ID>IN_1</ID>620 </input>
<input>
<ID>IN_2</ID>616 </input>
<input>
<ID>IN_3</ID>615 </input>
<output>
<ID>OUT</ID>623 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>472</ID>
<type>AE_OR2</type>
<position>437,1955.5</position>
<input>
<ID>IN_0</ID>623 </input>
<input>
<ID>IN_1</ID>624 </input>
<output>
<ID>OUT</ID>738 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>475</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>461,1962</position>
<input>
<ID>IN_0</ID>716 </input>
<input>
<ID>IN_1</ID>717 </input>
<input>
<ID>IN_2</ID>718 </input>
<input>
<ID>IN_3</ID>719 </input>
<output>
<ID>carry_out</ID>700 </output>
<input>
<ID>clear</ID>744 </input>
<input>
<ID>clock</ID>741 </input>
<input>
<ID>load</ID>598 </input>
<input>
<ID>shift_enable</ID>701 </input>
<input>
<ID>shift_left</ID>720 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>476</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>461,1949</position>
<input>
<ID>carry_in</ID>700 </input>
<input>
<ID>clear</ID>744 </input>
<input>
<ID>clock</ID>741 </input>
<input>
<ID>shift_enable</ID>701 </input>
<input>
<ID>shift_left</ID>739 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>477</ID>
<type>BB_CLOCK</type>
<position>406,1939</position>
<output>
<ID>CLK</ID>709 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>478</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>414,1945.5</position>
<input>
<ID>IN_0</ID>710 </input>
<output>
<ID>OUT_0</ID>711 </output>
<output>
<ID>OUT_1</ID>712 </output>
<output>
<ID>OUT_2</ID>713 </output>
<output>
<ID>OUT_3</ID>714 </output>
<output>
<ID>carry_out</ID>737 </output>
<input>
<ID>clear</ID>737 </input>
<input>
<ID>clock</ID>709 </input>
<input>
<ID>load</ID>738 </input>
<input>
<ID>shift_enable</ID>710 </input>
<input>
<ID>shift_left</ID>710 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>479</ID>
<type>EE_VDD</type>
<position>409.5,1947</position>
<output>
<ID>OUT_0</ID>710 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>480</ID>
<type>AE_OR4</type>
<position>422.5,1945.5</position>
<input>
<ID>IN_0</ID>711 </input>
<input>
<ID>IN_1</ID>712 </input>
<input>
<ID>IN_2</ID>713 </input>
<input>
<ID>IN_3</ID>714 </input>
<output>
<ID>OUT</ID>721 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>289</ID>
<type>AE_SMALL_INVERTER</type>
<position>451.5,1941.5</position>
<input>
<ID>IN_0</ID>599 </input>
<output>
<ID>OUT_0</ID>598 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>485</ID>
<type>GA_LED</type>
<position>435.5,1944.5</position>
<input>
<ID>N_in0</ID>735 </input>
<input>
<ID>N_in1</ID>715 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>AE_SMALL_INVERTER</type>
<position>439.5,1941.5</position>
<input>
<ID>IN_0</ID>601 </input>
<output>
<ID>OUT_0</ID>600 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>491</ID>
<type>DE_TO</type>
<position>438.5,1944.5</position>
<input>
<ID>IN_0</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cc</lparam></gate>
<gate>
<ID>492</ID>
<type>EE_VDD</type>
<position>463,1968</position>
<output>
<ID>OUT_0</ID>720 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>493</ID>
<type>EE_VDD</type>
<position>464,1956</position>
<output>
<ID>OUT_0</ID>739 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>494</ID>
<type>AA_AND2</type>
<position>431.5,1944.5</position>
<input>
<ID>IN_0</ID>721 </input>
<input>
<ID>IN_1</ID>736 </input>
<output>
<ID>OUT</ID>735 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>495</ID>
<type>AE_SMALL_INVERTER</type>
<position>418,1939</position>
<input>
<ID>IN_0</ID>709 </input>
<output>
<ID>OUT_0</ID>596 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>496</ID>
<type>AE_SMALL_INVERTER</type>
<position>422,1939</position>
<input>
<ID>IN_0</ID>596 </input>
<output>
<ID>OUT_0</ID>736 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>303</ID>
<type>AE_SMALL_INVERTER</type>
<position>443.5,1941.5</position>
<input>
<ID>IN_0</ID>600 </input>
<output>
<ID>OUT_0</ID>602 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>497</ID>
<type>DA_FROM</type>
<position>461,1973</position>
<input>
<ID>IN_0</ID>701 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID cc</lparam></gate>
<gate>
<ID>498</ID>
<type>AE_SMALL_INVERTER</type>
<position>439.5,1939</position>
<input>
<ID>IN_0</ID>736 </input>
<output>
<ID>OUT_0</ID>740 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>499</ID>
<type>AE_SMALL_INVERTER</type>
<position>443.5,1939</position>
<input>
<ID>IN_0</ID>740 </input>
<output>
<ID>OUT_0</ID>743 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>500</ID>
<type>AE_SMALL_INVERTER</type>
<position>447.5,1939</position>
<input>
<ID>IN_0</ID>743 </input>
<output>
<ID>OUT_0</ID>742 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>501</ID>
<type>AE_SMALL_INVERTER</type>
<position>451.5,1939</position>
<input>
<ID>IN_0</ID>742 </input>
<output>
<ID>OUT_0</ID>741 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>503</ID>
<type>CC_PULSE</type>
<position>399.5,1979.5</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>505</ID>
<type>CC_PULSE</type>
<position>399.5,1976.5</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>507</ID>
<type>CC_PULSE</type>
<position>399.5,1974</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>509</ID>
<type>CC_PULSE</type>
<position>399.5,1971.5</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>511</ID>
<type>CC_PULSE</type>
<position>399.5,1969</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>513</ID>
<type>CC_PULSE</type>
<position>399.5,1966.5</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>515</ID>
<type>CC_PULSE</type>
<position>399.5,1964</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>517</ID>
<type>CC_PULSE</type>
<position>399.5,1961</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>327</ID>
<type>DA_FROM</type>
<position>462,1929</position>
<input>
<ID>IN_0</ID>745 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>521</ID>
<type>DD_KEYPAD_HEX</type>
<position>491.5,1949.5</position>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>328</ID>
<type>DE_TO</type>
<position>447.5,1950</position>
<input>
<ID>IN_0</ID>738 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID klaw</lparam></gate>
<gate>
<ID>522</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>510.5,1967.5</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>166</ID>
<type>AE_SMALL_INVERTER</type>
<position>431.5,1941.5</position>
<input>
<ID>IN_0</ID>714 </input>
<output>
<ID>OUT_0</ID>597 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>167</ID>
<type>AE_SMALL_INVERTER</type>
<position>435.5,1941.5</position>
<input>
<ID>IN_0</ID>597 </input>
<output>
<ID>OUT_0</ID>601 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>168</ID>
<type>AE_SMALL_INVERTER</type>
<position>447.5,1941.5</position>
<input>
<ID>IN_0</ID>602 </input>
<output>
<ID>OUT_0</ID>599 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>560</ID>
<type>AE_REGISTER8</type>
<position>497.5,1962.5</position>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>420,1939,420,1939</points>
<connection>
<GID>495</GID>
<name>OUT_0</name></connection>
<connection>
<GID>496</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>433.5,1941.5,433.5,1941.5</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<connection>
<GID>167</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,1941.5,455.5,1969.5</points>
<intersection>1941.5 1</intersection>
<intersection>1969.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>453.5,1941.5,455.5,1941.5</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<intersection>455.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>455.5,1969.5,462,1969.5</points>
<intersection>455.5 0</intersection>
<intersection>462 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>462,1967,462,1969.5</points>
<connection>
<GID>475</GID>
<name>load</name></connection>
<intersection>1969.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449.5,1941.5,449.5,1941.5</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<connection>
<GID>289</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>441.5,1941.5,441.5,1941.5</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<connection>
<GID>303</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437.5,1941.5,437.5,1941.5</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<connection>
<GID>296</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445.5,1941.5,445.5,1941.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<connection>
<GID>303</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>412.5,1955.5,412.5,1963</points>
<intersection>1955.5 2</intersection>
<intersection>1963 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1963,412.5,1963</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>412.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>412.5,1955.5,419,1955.5</points>
<connection>
<GID>437</GID>
<name>IN_4</name></connection>
<intersection>412.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413,1956.5,413,1967</points>
<intersection>1956.5 2</intersection>
<intersection>1966 3</intersection>
<intersection>1967 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1967,413,1967</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413,1956.5,419,1956.5</points>
<connection>
<GID>437</GID>
<name>IN_5</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>413,1966,418,1966</points>
<connection>
<GID>440</GID>
<name>IN_2</name></connection>
<intersection>413 0</intersection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413.5,1957.5,413.5,1974</points>
<intersection>1957.5 2</intersection>
<intersection>1971 1</intersection>
<intersection>1974 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1971,413.5,1971</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>413.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413.5,1957.5,419,1957.5</points>
<connection>
<GID>437</GID>
<name>IN_6</name></connection>
<intersection>413.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>413.5,1974,418,1974</points>
<connection>
<GID>441</GID>
<name>IN_2</name></connection>
<intersection>413.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>414,1958.5,414,1978</points>
<intersection>1958.5 2</intersection>
<intersection>1970 3</intersection>
<intersection>1975 1</intersection>
<intersection>1978 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1975,414,1975</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>414 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>414,1958.5,419,1958.5</points>
<connection>
<GID>437</GID>
<name>IN_7</name></connection>
<intersection>414 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>414,1970,418,1970</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>414 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>414,1978,418,1978</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>414 0</intersection></hsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>414.5,1959.5,414.5,1982</points>
<intersection>1959.5 2</intersection>
<intersection>1979 1</intersection>
<intersection>1982 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1979,414.5,1979</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<intersection>414.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>414.5,1959.5,419,1959.5</points>
<connection>
<GID>437</GID>
<name>IN_3</name></connection>
<intersection>414.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>414.5,1982,419,1982</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<intersection>414.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>419,1960.5,419,1962.5</points>
<connection>
<GID>438</GID>
<name>OUT_0</name></connection>
<connection>
<GID>437</GID>
<name>IN_2</name></connection>
<connection>
<GID>437</GID>
<name>IN_1</name></connection>
<connection>
<GID>437</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426,1956,426,1969</points>
<connection>
<GID>437</GID>
<name>OUT</name></connection>
<intersection>1956 6</intersection>
<intersection>1969 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>426,1969,430,1969</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<intersection>426 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>426,1956,427,1956</points>
<connection>
<GID>471</GID>
<name>IN_3</name></connection>
<intersection>426 0</intersection></hsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,1958,425.5,1970</points>
<intersection>1958 3</intersection>
<intersection>1967 2</intersection>
<intersection>1970 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425.5,1970,430,1970</points>
<connection>
<GID>436</GID>
<name>IN_1</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>425,1967,425.5,1967</points>
<connection>
<GID>440</GID>
<name>OUT</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>425.5,1958,427,1958</points>
<connection>
<GID>471</GID>
<name>IN_2</name></connection>
<intersection>425.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413,1964,413,1965</points>
<intersection>1964 2</intersection>
<intersection>1965 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1965,413,1965</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413,1964,418,1964</points>
<connection>
<GID>440</GID>
<name>IN_3</name></connection>
<intersection>413 0</intersection></hsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413,1968,413,1976</points>
<intersection>1968 2</intersection>
<intersection>1973 1</intersection>
<intersection>1976 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1973,413,1973</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413,1968,418,1968</points>
<connection>
<GID>440</GID>
<name>IN_1</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>413,1976,418,1976</points>
<connection>
<GID>441</GID>
<name>IN_1</name></connection>
<intersection>413 0</intersection></hsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426,1972,426,1981</points>
<intersection>1972 3</intersection>
<intersection>1981 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>425,1981,426,1981</points>
<connection>
<GID>439</GID>
<name>OUT</name></connection>
<intersection>426 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>426,1972,430,1972</points>
<connection>
<GID>436</GID>
<name>IN_3</name></connection>
<intersection>426 0</intersection>
<intersection>427 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>427,1962,427,1972</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<intersection>1972 3</intersection></vsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,1971,425.5,1975</points>
<intersection>1971 1</intersection>
<intersection>1975 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425.5,1971,430,1971</points>
<connection>
<GID>436</GID>
<name>IN_2</name></connection>
<intersection>425.5 0</intersection>
<intersection>426.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>425,1975,425.5,1975</points>
<connection>
<GID>441</GID>
<name>OUT</name></connection>
<intersection>425.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>426.5,1960,426.5,1971</points>
<intersection>1960 6</intersection>
<intersection>1971 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>426.5,1960,427,1960</points>
<connection>
<GID>471</GID>
<name>IN_1</name></connection>
<intersection>426.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413.5,1977,413.5,1980</points>
<intersection>1977 1</intersection>
<intersection>1980 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1977,413.5,1977</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<intersection>413.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413.5,1980,419,1980</points>
<connection>
<GID>439</GID>
<name>IN_1</name></connection>
<intersection>413.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413,1969,413,1972</points>
<intersection>1969 1</intersection>
<intersection>1972 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1969,413,1969</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413,1972,418,1972</points>
<connection>
<GID>441</GID>
<name>IN_3</name></connection>
<intersection>413 0</intersection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>434,1956.5,434,1959</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<connection>
<GID>471</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>412,1954.5,412,1961</points>
<intersection>1954.5 2</intersection>
<intersection>1961 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1961,412,1961</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>412 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>412,1954.5,434,1954.5</points>
<connection>
<GID>472</GID>
<name>IN_1</name></connection>
<intersection>412 0</intersection></hsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431.5,1962.5,431.5,1966</points>
<connection>
<GID>436</GID>
<name>OUT_3</name></connection>
<intersection>1962.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>431.5,1962.5,437,1962.5</points>
<connection>
<GID>433</GID>
<name>IN_3</name></connection>
<intersection>431.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432.5,1961.5,432.5,1966</points>
<connection>
<GID>436</GID>
<name>OUT_2</name></connection>
<intersection>1961.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,1961.5,437,1961.5</points>
<connection>
<GID>433</GID>
<name>IN_2</name></connection>
<intersection>432.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>433.5,1960.5,433.5,1966</points>
<connection>
<GID>436</GID>
<name>OUT_1</name></connection>
<intersection>1960.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>433.5,1960.5,437,1960.5</points>
<connection>
<GID>433</GID>
<name>IN_1</name></connection>
<intersection>433.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,1959.5,434.5,1966</points>
<connection>
<GID>436</GID>
<name>OUT_0</name></connection>
<intersection>1959.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,1959.5,437,1959.5</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<vsegment>
<ID>20</ID>
<points>459.5,1954,459.5,1957</points>
<connection>
<GID>476</GID>
<name>carry_in</name></connection>
<connection>
<GID>475</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>466,1954.5,466,1971</points>
<intersection>1954.5 20</intersection>
<intersection>1971 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>461,1971,466,1971</points>
<intersection>461 22</intersection>
<intersection>466 1</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>461,1954.5,466,1954.5</points>
<intersection>461 21</intersection>
<intersection>466 1</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>461,1954,461,1954.5</points>
<connection>
<GID>476</GID>
<name>shift_enable</name></connection>
<intersection>1954.5 20</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>461,1967,461,1971</points>
<connection>
<GID>475</GID>
<name>shift_enable</name></connection>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<intersection>1971 18</intersection></vsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<vsegment>
<ID>18</ID>
<points>415,1939,415,1940.5</points>
<connection>
<GID>478</GID>
<name>clock</name></connection>
<intersection>1939 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>410,1939,416,1939</points>
<connection>
<GID>477</GID>
<name>CLK</name></connection>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>415 18</intersection></hsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>410.5,1947,410.5,1951.5</points>
<connection>
<GID>479</GID>
<name>OUT_0</name></connection>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>1951.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>410.5,1951.5,416,1951.5</points>
<intersection>410.5 0</intersection>
<intersection>414 14</intersection>
<intersection>416 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>416,1950.5,416,1951.5</points>
<connection>
<GID>478</GID>
<name>shift_left</name></connection>
<intersection>1951.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>414,1950.5,414,1951.5</points>
<connection>
<GID>478</GID>
<name>shift_enable</name></connection>
<intersection>1951.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>418,1947,418,1948.5</points>
<intersection>1947 1</intersection>
<intersection>1948.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>417.5,1947,418,1947</points>
<connection>
<GID>478</GID>
<name>OUT_0</name></connection>
<intersection>418 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>418,1948.5,419.5,1948.5</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>418 0</intersection></hsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>417.5,1946.5,419.5,1946.5</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>417.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>417.5,1946,417.5,1946.5</points>
<connection>
<GID>478</GID>
<name>OUT_1</name></connection>
<intersection>1946.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>417.5,1944.5,419.5,1944.5</points>
<connection>
<GID>480</GID>
<name>IN_2</name></connection>
<intersection>417.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>417.5,1944.5,417.5,1945</points>
<connection>
<GID>478</GID>
<name>OUT_2</name></connection>
<intersection>1944.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>417.5,1941.5,417.5,1944</points>
<connection>
<GID>478</GID>
<name>OUT_3</name></connection>
<intersection>1941.5 12</intersection>
<intersection>1942.5 15</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>417.5,1941.5,429.5,1941.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>417.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>417.5,1942.5,419.5,1942.5</points>
<connection>
<GID>480</GID>
<name>IN_3</name></connection>
<intersection>417.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436.5,1944.5,436.5,1944.5</points>
<connection>
<GID>485</GID>
<name>N_in1</name></connection>
<connection>
<GID>491</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>453,1959.5,453,1963.5</points>
<intersection>1959.5 1</intersection>
<intersection>1963.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445,1959.5,453,1959.5</points>
<connection>
<GID>433</GID>
<name>OUT_0</name></connection>
<intersection>453 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>453,1963.5,457.5,1963.5</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>453 0</intersection></hsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448.5,1960.5,448.5,1963</points>
<intersection>1960.5 1</intersection>
<intersection>1963 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445,1960.5,448.5,1960.5</points>
<connection>
<GID>433</GID>
<name>OUT_1</name></connection>
<intersection>448.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448.5,1963,457.5,1963</points>
<intersection>448.5 0</intersection>
<intersection>457.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>457.5,1962.5,457.5,1963</points>
<connection>
<GID>475</GID>
<name>IN_1</name></connection>
<intersection>1963 2</intersection></vsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>445,1961.5,457.5,1961.5</points>
<connection>
<GID>433</GID>
<name>OUT_2</name></connection>
<connection>
<GID>475</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450,1960.5,450,1962.5</points>
<intersection>1960.5 2</intersection>
<intersection>1962.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445,1962.5,450,1962.5</points>
<connection>
<GID>433</GID>
<name>OUT_3</name></connection>
<intersection>450 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450,1960.5,457.5,1960.5</points>
<connection>
<GID>475</GID>
<name>IN_3</name></connection>
<intersection>450 0</intersection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>463,1967,463,1967</points>
<connection>
<GID>475</GID>
<name>shift_left</name></connection>
<connection>
<GID>492</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>426.5,1945.5,428.5,1945.5</points>
<connection>
<GID>480</GID>
<name>OUT</name></connection>
<connection>
<GID>494</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,1944.5,434.5,1944.5</points>
<connection>
<GID>485</GID>
<name>N_in0</name></connection>
<connection>
<GID>494</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428,1939,428,1943.5</points>
<intersection>1939 5</intersection>
<intersection>1943.5 15</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>424,1939,437.5,1939</points>
<connection>
<GID>496</GID>
<name>OUT_0</name></connection>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>428 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>428,1943.5,428.5,1943.5</points>
<connection>
<GID>494</GID>
<name>IN_1</name></connection>
<intersection>428 0</intersection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412.5,1940.5,414,1940.5</points>
<connection>
<GID>478</GID>
<name>clear</name></connection>
<connection>
<GID>478</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>415,1950.5,415,1953</points>
<connection>
<GID>478</GID>
<name>load</name></connection>
<intersection>1953 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>415,1953,447,1953</points>
<intersection>415 0</intersection>
<intersection>445.5 16</intersection>
<intersection>447 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>447,1953,447,1973</points>
<intersection>1953 1</intersection>
<intersection>1955.5 5</intersection>
<intersection>1973 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>440,1973,447,1973</points>
<intersection>440 7</intersection>
<intersection>447 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>440,1955.5,447,1955.5</points>
<connection>
<GID>472</GID>
<name>OUT</name></connection>
<intersection>440 8</intersection>
<intersection>447 2</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>440,1968.5,440,1973</points>
<connection>
<GID>433</GID>
<name>load</name></connection>
<intersection>1973 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>440,1955.5,440,1957.5</points>
<connection>
<GID>433</GID>
<name>clock</name></connection>
<intersection>1955.5 5</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>445.5,1950,445.5,1953</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>1953 1</intersection></vsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>463,1954,463,1956</points>
<connection>
<GID>493</GID>
<name>OUT_0</name></connection>
<connection>
<GID>476</GID>
<name>shift_left</name></connection></vsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>441.5,1939,441.5,1939</points>
<connection>
<GID>498</GID>
<name>OUT_0</name></connection>
<connection>
<GID>499</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>465,1939,465,1957</points>
<intersection>1939 8</intersection>
<intersection>1944 5</intersection>
<intersection>1957 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>462,1944,465,1944</points>
<connection>
<GID>476</GID>
<name>clock</name></connection>
<intersection>465 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>462,1957,465,1957</points>
<connection>
<GID>475</GID>
<name>clock</name></connection>
<intersection>465 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>453.5,1939,465,1939</points>
<connection>
<GID>501</GID>
<name>OUT_0</name></connection>
<intersection>465 0</intersection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449.5,1939,449.5,1939</points>
<connection>
<GID>500</GID>
<name>OUT_0</name></connection>
<connection>
<GID>501</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445.5,1939,445.5,1939</points>
<connection>
<GID>499</GID>
<name>OUT_0</name></connection>
<connection>
<GID>500</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>744</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454.5,1940,454.5,1957</points>
<intersection>1940 4</intersection>
<intersection>1957 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>454.5,1957,461,1957</points>
<connection>
<GID>475</GID>
<name>clear</name></connection>
<intersection>454.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>454.5,1940,461,1940</points>
<intersection>454.5 0</intersection>
<intersection>461 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>461,1937,461,1944</points>
<connection>
<GID>434</GID>
<name>OUT</name></connection>
<connection>
<GID>476</GID>
<name>clear</name></connection>
<intersection>1940 4</intersection></vsegment></shape></wire>
<wire>
<ID>745</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>462,1931,462,1931</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<connection>
<GID>434</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>746</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>460,1931,460,1931</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<connection>
<GID>435</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-22.5313,2284.15,1755.47,1357.15</PageViewport></page 5>
<page 6>
<PageViewport>-22.5313,2284.15,1755.47,1357.15</PageViewport></page 6>
<page 7>
<PageViewport>-22.5313,2284.15,1755.47,1357.15</PageViewport></page 7>
<page 8>
<PageViewport>-22.5313,2284.15,1755.47,1357.15</PageViewport></page 8>
<page 9>
<PageViewport>-22.5313,2284.15,1755.47,1357.15</PageViewport></page 9></circuit>