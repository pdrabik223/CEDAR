<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>24.6333,-8.33333,261.7,-131.933</PageViewport>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>84.5,-22.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_DFF_LOW</type>
<position>127,-24</position>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>32</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>65,-15</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>34</ID>
<type>BE_JKFF_LOW</type>
<position>103.5,-35</position>
<input>
<ID>J</ID>5 </input>
<input>
<ID>K</ID>5 </input>
<output>
<ID>Q</ID>24 </output>
<input>
<ID>clock</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>46</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>58.5,-15</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>47</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>52,-15</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>56</ID>
<type>GA_LED</type>
<position>36.5,-14.5</position>
<input>
<ID>N_in0</ID>23 </input>
<input>
<ID>N_in1</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>GA_LED</type>
<position>38.5,-14.5</position>
<input>
<ID>N_in0</ID>22 </input>
<input>
<ID>N_in1</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>40.5,-14.5</position>
<input>
<ID>N_in0</ID>22 </input>
<input>
<ID>N_in1</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>42.5,-14.5</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>DA_FROM</type>
<position>33.5,-14.5</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID om</lparam></gate>
<gate>
<ID>65</ID>
<type>DE_TO</type>
<position>108.5,-33</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID om</lparam></gate>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>86.5,-35,100.5,-35</points>
<connection>
<GID>34</GID>
<name>clock</name></connection>
<intersection>86.5 3</intersection>
<intersection>100.5 18</intersection>
<intersection>100.5 18</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>86.5,-35,86.5,-22.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-35 2</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>100.5,-37,100.5,-33</points>
<connection>
<GID>34</GID>
<name>J</name></connection>
<connection>
<GID>34</GID>
<name>K</name></connection>
<intersection>-35 2</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>41.5,-14.5,41.5,-14.5</points>
<connection>
<GID>58</GID>
<name>N_in1</name></connection>
<connection>
<GID>59</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-14.5,39.5,-14.5</points>
<connection>
<GID>56</GID>
<name>N_in1</name></connection>
<connection>
<GID>57</GID>
<name>N_in0</name></connection>
<connection>
<GID>57</GID>
<name>N_in1</name></connection>
<connection>
<GID>58</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-14.5,35.5,-14.5</points>
<connection>
<GID>56</GID>
<name>N_in0</name></connection>
<connection>
<GID>60</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-33,106.5,-33</points>
<connection>
<GID>34</GID>
<name>Q</name></connection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-33,106.5,-33</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>4.36481,19.4949,122.898,-42.3051</PageViewport>
<gate>
<ID>194</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>99.5,-4</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>176 </input>
<input>
<ID>IN_2</ID>177 </input>
<input>
<ID>IN_3</ID>178 </input>
<output>
<ID>OUT_0</ID>198 </output>
<output>
<ID>OUT_1</ID>197 </output>
<output>
<ID>OUT_2</ID>196 </output>
<output>
<ID>OUT_3</ID>195 </output>
<output>
<ID>carry_out</ID>120 </output>
<input>
<ID>clear</ID>180 </input>
<input>
<ID>clock</ID>121 </input>
<input>
<ID>shift_enable</ID>122 </input>
<input>
<ID>shift_left</ID>181 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>196</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>116,-10</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>197 </input>
<input>
<ID>IN_2</ID>196 </input>
<input>
<ID>IN_3</ID>195 </input>
<input>
<ID>IN_4</ID>194 </input>
<input>
<ID>IN_5</ID>193 </input>
<input>
<ID>IN_6</ID>192 </input>
<input>
<ID>IN_7</ID>191 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 144</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>197</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>99.5,-15</position>
<output>
<ID>OUT_0</ID>194 </output>
<output>
<ID>OUT_1</ID>193 </output>
<output>
<ID>OUT_2</ID>192 </output>
<output>
<ID>OUT_3</ID>191 </output>
<input>
<ID>carry_in</ID>120 </input>
<input>
<ID>clear</ID>180 </input>
<input>
<ID>clock</ID>121 </input>
<input>
<ID>shift_enable</ID>179 </input>
<input>
<ID>shift_left</ID>182 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>201</ID>
<type>CC_PULSE</type>
<position>15,0</position>
<output>
<ID>OUT_0</ID>226 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 9</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>205</ID>
<type>BB_CLOCK</type>
<position>35,-28.5</position>
<output>
<ID>CLK</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>237</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>47,-22</position>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUT_0</ID>167 </output>
<output>
<ID>OUT_1</ID>168 </output>
<output>
<ID>OUT_2</ID>169 </output>
<output>
<ID>OUT_3</ID>170 </output>
<output>
<ID>carry_out</ID>220 </output>
<input>
<ID>clear</ID>220 </input>
<input>
<ID>clock</ID>152 </input>
<input>
<ID>load</ID>225 </input>
<input>
<ID>shift_enable</ID>160 </input>
<input>
<ID>shift_left</ID>160 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>239</ID>
<type>EE_VDD</type>
<position>42,-19.5</position>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>243</ID>
<type>AE_OR4</type>
<position>55.5,-22</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>168 </input>
<input>
<ID>IN_2</ID>169 </input>
<input>
<ID>IN_3</ID>170 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>247</ID>
<type>GA_LED</type>
<position>66.5,-23</position>
<input>
<ID>N_in0</ID>206 </input>
<input>
<ID>N_in1</ID>174 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>249</ID>
<type>DE_TO</type>
<position>69.5,-23</position>
<input>
<ID>IN_0</ID>174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cc</lparam></gate>
<gate>
<ID>250</ID>
<type>BB_CLOCK</type>
<position>92.5,-25</position>
<output>
<ID>CLK</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_AND2</type>
<position>106,7</position>
<input>
<ID>IN_0</ID>122 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>CC_PULSE</type>
<position>86.5,-21.5</position>
<output>
<ID>OUT_0</ID>180 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 9</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>255</ID>
<type>EE_VDD</type>
<position>101.5,2.5</position>
<output>
<ID>OUT_0</ID>181 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>256</ID>
<type>EE_VDD</type>
<position>107.5,-10</position>
<output>
<ID>OUT_0</ID>182 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>262</ID>
<type>DE_TO</type>
<position>39,-33</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID TO</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_AND2</type>
<position>62.5,-23</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>218 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>269</ID>
<type>AE_SMALL_INVERTER</type>
<position>50,-28.5</position>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT_0</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>270</ID>
<type>AE_SMALL_INVERTER</type>
<position>54,-28.5</position>
<input>
<ID>IN_0</ID>213 </input>
<output>
<ID>OUT_0</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>278</ID>
<type>DA_FROM</type>
<position>100,13</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID cc</lparam></gate>
<gate>
<ID>280</ID>
<type>DE_TO</type>
<position>19,0</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID load</lparam></gate>
<gate>
<ID>284</ID>
<type>DA_FROM</type>
<position>95.5,6.5</position>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID load</lparam></gate>
<gate>
<ID>285</ID>
<type>DA_FROM</type>
<position>25.5,-17</position>
<input>
<ID>IN_0</ID>224 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID load</lparam></gate>
<gate>
<ID>286</ID>
<type>AE_SMALL_INVERTER</type>
<position>29.5,-17</position>
<input>
<ID>IN_0</ID>224 </input>
<output>
<ID>OUT_0</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>287</ID>
<type>AE_SMALL_INVERTER</type>
<position>33.5,-17</position>
<input>
<ID>IN_0</ID>223 </input>
<output>
<ID>OUT_0</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>96</ID>
<type>DA_FROM</type>
<position>45,-2</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>97</ID>
<type>DA_FROM</type>
<position>45,0</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>98</ID>
<type>DA_FROM</type>
<position>45,2</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>99</ID>
<type>DA_FROM</type>
<position>45,4</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>45,6</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>45,8</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>45,10</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>103</ID>
<type>DA_FROM</type>
<position>45,12</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>104</ID>
<type>DA_FROM</type>
<position>45,14</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>107</ID>
<type>AE_REGISTER8</type>
<position>79.5,-2.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>109 </input>
<input>
<ID>IN_2</ID>108 </input>
<input>
<ID>IN_3</ID>107 </input>
<output>
<ID>OUT_0</ID>175 </output>
<output>
<ID>OUT_1</ID>176 </output>
<output>
<ID>OUT_2</ID>177 </output>
<output>
<ID>OUT_3</ID>178 </output>
<input>
<ID>clock</ID>106 </input>
<input>
<ID>load</ID>106 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 8</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>117</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-23,5</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>119</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>71.5,5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>78 </input>
<input>
<ID>IN_2</ID>82 </input>
<input>
<ID>IN_3</ID>81 </input>
<output>
<ID>OUT_0</ID>110 </output>
<output>
<ID>OUT_1</ID>109 </output>
<output>
<ID>OUT_2</ID>108 </output>
<output>
<ID>OUT_3</ID>107 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>134</ID>
<type>BA_DECODER_2x4</type>
<position>4,-2</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_OR8</type>
<position>60.5,-6</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>69 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>68 </input>
<input>
<ID>IN_4</ID>64 </input>
<input>
<ID>IN_5</ID>65 </input>
<input>
<ID>IN_6</ID>66 </input>
<input>
<ID>IN_7</ID>67 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>140</ID>
<type>FF_GND</type>
<position>56.5,-4.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>145</ID>
<type>AE_OR2</type>
<position>60.5,16</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_OR4</type>
<position>59.5,2</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>80 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>79 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>148</ID>
<type>AE_OR4</type>
<position>59.5,10</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>80 </input>
<input>
<ID>IN_2</ID>66 </input>
<input>
<ID>IN_3</ID>84 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>149</ID>
<type>CC_PULSE</type>
<position>32,-13.5</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>150</ID>
<type>CC_PULSE</type>
<position>36,9</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>151</ID>
<type>CC_PULSE</type>
<position>32,9</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>152</ID>
<type>CC_PULSE</type>
<position>28,9</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>153</ID>
<type>CC_PULSE</type>
<position>36,1.5</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>154</ID>
<type>CC_PULSE</type>
<position>32,1.5</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>155</ID>
<type>CC_PULSE</type>
<position>28,1.5</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>156</ID>
<type>CC_PULSE</type>
<position>36,-6</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>157</ID>
<type>CC_PULSE</type>
<position>32,-6</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>158</ID>
<type>CC_PULSE</type>
<position>28,-6</position>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>159</ID>
<type>DE_TO</type>
<position>28,13</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>160</ID>
<type>DE_TO</type>
<position>32,13</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>161</ID>
<type>DE_TO</type>
<position>36,13</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>162</ID>
<type>DE_TO</type>
<position>28,5.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>163</ID>
<type>DE_TO</type>
<position>32,5.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>164</ID>
<type>DE_TO</type>
<position>36,5.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>165</ID>
<type>DE_TO</type>
<position>28,-2</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>166</ID>
<type>DE_TO</type>
<position>32,-2</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>167</ID>
<type>DE_TO</type>
<position>36,-2</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_TO</type>
<position>32,-9.5</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>172</ID>
<type>GA_LED</type>
<position>10.5,2</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>45,-4</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>183</ID>
<type>AE_OR4</type>
<position>68.5,-6</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>78 </input>
<input>
<ID>IN_3</ID>77 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>185</ID>
<type>AE_OR2</type>
<position>75.5,-9.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-14.5,107,-8</points>
<intersection>-14.5 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-8,111,-8</points>
<connection>
<GID>196</GID>
<name>IN_5</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-14.5,107,-14.5</points>
<connection>
<GID>197</GID>
<name>OUT_1</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-13.5,107,-9</points>
<intersection>-13.5 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-9,111,-9</points>
<connection>
<GID>196</GID>
<name>IN_4</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-13.5,107,-13.5</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-10,107,-5.5</points>
<intersection>-10 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-10,111,-10</points>
<connection>
<GID>196</GID>
<name>IN_3</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-5.5,107,-5.5</points>
<connection>
<GID>194</GID>
<name>OUT_3</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-11,107,-4.5</points>
<intersection>-11 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-11,111,-11</points>
<connection>
<GID>196</GID>
<name>IN_2</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-4.5,107,-4.5</points>
<connection>
<GID>194</GID>
<name>OUT_2</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-12,107,-3.5</points>
<intersection>-12 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-12,111,-12</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-3.5,107,-3.5</points>
<connection>
<GID>194</GID>
<name>OUT_1</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-13,107,-2.5</points>
<intersection>-13 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-13,111,-13</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-2.5,107,-2.5</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-22,59.5,-22</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<connection>
<GID>263</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-23,65.5,-23</points>
<connection>
<GID>247</GID>
<name>N_in0</name></connection>
<connection>
<GID>263</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-28.5,52,-28.5</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-28.5,59.5,-24</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<intersection>-28.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>56,-28.5,59.5,-28.5</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-27,47,-27</points>
<connection>
<GID>237</GID>
<name>clear</name></connection>
<connection>
<GID>237</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-17,31.5,-17</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-17,27.5,-17</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<connection>
<GID>286</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-14.5,48,-14.5</points>
<intersection>35.5 3</intersection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-17,48,-14.5</points>
<connection>
<GID>237</GID>
<name>load</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-17,35.5,-14.5</points>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,0,17,0</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-9.5,51,-2</points>
<intersection>-9.5 2</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-2,51,-2</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-9.5,57.5,-9.5</points>
<connection>
<GID>138</GID>
<name>IN_4</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-8.5,51.5,2</points>
<intersection>-8.5 2</intersection>
<intersection>1 3</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,2,51.5,2</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-8.5,57.5,-8.5</points>
<connection>
<GID>138</GID>
<name>IN_5</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51.5,1,56.5,1</points>
<connection>
<GID>147</GID>
<name>IN_2</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-7.5,52,9</points>
<intersection>-7.5 2</intersection>
<intersection>6 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,6,52,6</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-7.5,57.5,-7.5</points>
<connection>
<GID>138</GID>
<name>IN_6</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52,9,56.5,9</points>
<connection>
<GID>148</GID>
<name>IN_2</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-6.5,52.5,13</points>
<intersection>-6.5 2</intersection>
<intersection>5 3</intersection>
<intersection>10 1</intersection>
<intersection>13 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,10,52.5,10</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-6.5,57.5,-6.5</points>
<connection>
<GID>138</GID>
<name>IN_7</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52.5,5,56.5,5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,13,56.5,13</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-5.5,53,17</points>
<intersection>-5.5 2</intersection>
<intersection>14 1</intersection>
<intersection>17 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,14,53,14</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-5.5,57.5,-5.5</points>
<connection>
<GID>138</GID>
<name>IN_3</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>53,17,57.5,17</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-4.5,57.5,-2.5</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<connection>
<GID>138</GID>
<name>IN_2</name></connection>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-9,64.5,4</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>-9 6</intersection>
<intersection>4 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>64.5,4,68.5,4</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>64.5,-9,65.5,-9</points>
<connection>
<GID>183</GID>
<name>IN_3</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-7,64,5</points>
<intersection>-7 3</intersection>
<intersection>2 2</intersection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,5,68.5,5</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,2,64,2</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,-7,65.5,-7</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-1,51.5,0</points>
<intersection>-1 2</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,0,51.5,0</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-1,56.5,-1</points>
<connection>
<GID>147</GID>
<name>IN_3</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,3,51.5,11</points>
<intersection>3 2</intersection>
<intersection>8 1</intersection>
<intersection>11 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,8,51.5,8</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,3,56.5,3</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51.5,11,56.5,11</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,7,64.5,16</points>
<intersection>7 3</intersection>
<intersection>16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63.5,16,64.5,16</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64.5,7,68.5,7</points>
<connection>
<GID>119</GID>
<name>IN_3</name></connection>
<intersection>64.5 0</intersection>
<intersection>65.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>65.5,-3,65.5,7</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>7 3</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,6,64,10</points>
<intersection>6 1</intersection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,6,68.5,6</points>
<connection>
<GID>119</GID>
<name>IN_2</name></connection>
<intersection>64 0</intersection>
<intersection>65 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,10,64,10</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>64 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>65,-5,65,6</points>
<intersection>-5 6</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>65,-5,65.5,-5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>65 5</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,12,52,15</points>
<intersection>12 1</intersection>
<intersection>15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,12,52,12</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,15,57.5,15</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,4,51.5,7</points>
<intersection>4 1</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,4,51.5,4</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,7,56.5,7</points>
<connection>
<GID>148</GID>
<name>IN_3</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,11,28,11</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,11,28,11</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,11,32,11</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,11,36,11</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,3.5,28,3.5</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,3.5,32,3.5</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<connection>
<GID>163</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>36,3.5,36,3.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<connection>
<GID>164</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-4,28,-4</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<connection>
<GID>165</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-4,32,-4</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<connection>
<GID>166</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-4,36,-4</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<connection>
<GID>167</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-11.5,32,-11.5</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<connection>
<GID>168</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>72.5,-8.5,72.5,-6</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<connection>
<GID>185</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-10.5,50.5,-4</points>
<intersection>-10.5 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-4,50.5,-4</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-10.5,72.5,-10.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-9.5,89.5,5.5</points>
<intersection>-9.5 1</intersection>
<intersection>5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-9.5,89.5,-9.5</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>78.5 4</intersection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78.5,5.5,89.5,5.5</points>
<intersection>78.5 3</intersection>
<intersection>89.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>78.5,3.5,78.5,5.5</points>
<connection>
<GID>107</GID>
<name>load</name></connection>
<intersection>5.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-9.5,78.5,-7.5</points>
<connection>
<GID>107</GID>
<name>clock</name></connection>
<intersection>-9.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-2.5,70,1</points>
<connection>
<GID>119</GID>
<name>OUT_3</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-2.5,75.5,-2.5</points>
<connection>
<GID>107</GID>
<name>IN_3</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-3.5,71,1</points>
<connection>
<GID>119</GID>
<name>OUT_2</name></connection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-3.5,75.5,-3.5</points>
<connection>
<GID>107</GID>
<name>IN_2</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-4.5,72,1</points>
<connection>
<GID>119</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-4.5,75.5,-4.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-5.5,73,1</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-5.5,75.5,-5.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-10,98,-9</points>
<connection>
<GID>194</GID>
<name>carry_out</name></connection>
<connection>
<GID>197</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-27.5,105,-9</points>
<intersection>-27.5 4</intersection>
<intersection>-9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100.5,-9,105,-9</points>
<connection>
<GID>194</GID>
<name>clock</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>100.5,-27.5,105,-27.5</points>
<intersection>100.5 6</intersection>
<intersection>105 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>100.5,-27.5,100.5,-20</points>
<connection>
<GID>197</GID>
<name>clock</name></connection>
<intersection>-27.5 4</intersection>
<intersection>-25 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>96.5,-25,100.5,-25</points>
<connection>
<GID>250</GID>
<name>CLK</name></connection>
<intersection>100.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>100,6,100,11</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>6 2</intersection>
<intersection>10 8</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>99.5,6,100,6</points>
<intersection>99.5 6</intersection>
<intersection>100 1</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>99.5,1,99.5,6</points>
<connection>
<GID>194</GID>
<name>shift_enable</name></connection>
<intersection>6 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>100,10,107,10</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<connection>
<GID>251</GID>
<name>IN_1</name></connection>
<intersection>100 1</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>39,-28.5,48,-28.5</points>
<connection>
<GID>205</GID>
<name>CLK</name></connection>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>39 22</intersection>
<intersection>48 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>48,-28.5,48,-27</points>
<connection>
<GID>237</GID>
<name>clock</name></connection>
<intersection>-28.5 3</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>39,-31,39,-28.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>-28.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-20.5,43,-16.5</points>
<intersection>-20.5 1</intersection>
<intersection>-20 10</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-20.5,43.5,-20.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-16.5,49,-16.5</points>
<intersection>43 0</intersection>
<intersection>47 14</intersection>
<intersection>49 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>49,-17,49,-16.5</points>
<connection>
<GID>237</GID>
<name>shift_left</name></connection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>42.5,-20,43,-20</points>
<intersection>42.5 11</intersection>
<intersection>43 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>42.5,-20.5,42.5,-20</points>
<intersection>-20.5 12</intersection>
<intersection>-20 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>42,-20.5,42.5,-20.5</points>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection>
<intersection>42.5 11</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>47,-17,47,-16.5</points>
<connection>
<GID>237</GID>
<name>shift_enable</name></connection>
<intersection>-16.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-20.5,51,-19</points>
<intersection>-20.5 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-20.5,51,-20.5</points>
<connection>
<GID>237</GID>
<name>OUT_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-19,52.5,-19</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-21.5,52.5,-21.5</points>
<connection>
<GID>237</GID>
<name>OUT_1</name></connection>
<intersection>52.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>52.5,-21.5,52.5,-21</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>-21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-22.5,52.5,-22.5</points>
<connection>
<GID>237</GID>
<name>OUT_2</name></connection>
<intersection>52.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>52.5,-23,52.5,-22.5</points>
<connection>
<GID>243</GID>
<name>IN_2</name></connection>
<intersection>-22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-25,50.5,-23.5</points>
<connection>
<GID>237</GID>
<name>OUT_3</name></connection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-25,52.5,-25</points>
<connection>
<GID>243</GID>
<name>IN_3</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-23,67.5,-23</points>
<connection>
<GID>247</GID>
<name>N_in1</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-23,67.5,-23</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-5.5,89.5,-2.5</points>
<intersection>-5.5 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-5.5,89.5,-5.5</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-2.5,96,-2.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-4.5,89.5,-3.5</points>
<intersection>-4.5 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-4.5,89.5,-4.5</points>
<connection>
<GID>107</GID>
<name>OUT_1</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-3.5,96,-3.5</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-4.5,89.5,-3.5</points>
<intersection>-4.5 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-3.5,89.5,-3.5</points>
<connection>
<GID>107</GID>
<name>OUT_2</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-4.5,96,-4.5</points>
<connection>
<GID>194</GID>
<name>IN_2</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-5.5,89.5,-2.5</points>
<intersection>-5.5 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-2.5,89.5,-2.5</points>
<connection>
<GID>107</GID>
<name>OUT_3</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-5.5,96,-5.5</points>
<connection>
<GID>194</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-9.5,104.5,4</points>
<intersection>-9.5 2</intersection>
<intersection>4 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>99.5,-10,99.5,-9.5</points>
<connection>
<GID>197</GID>
<name>shift_enable</name></connection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>99.5,-9.5,104.5,-9.5</points>
<intersection>99.5 1</intersection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,4,106,4</points>
<connection>
<GID>251</GID>
<name>OUT</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-21.5,90.5,-9.5</points>
<intersection>-21.5 1</intersection>
<intersection>-20 4</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-21.5,90.5,-21.5</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>90.5,-9.5,99.5,-9.5</points>
<intersection>90.5 0</intersection>
<intersection>99.5 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>90.5,-20,99.5,-20</points>
<connection>
<GID>197</GID>
<name>clear</name></connection>
<intersection>90.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>99.5,-9.5,99.5,-9</points>
<connection>
<GID>194</GID>
<name>clear</name></connection>
<intersection>-9.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,1,101.5,1.5</points>
<connection>
<GID>194</GID>
<name>shift_left</name></connection>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101.5,-10,106.5,-10</points>
<connection>
<GID>197</GID>
<name>shift_left</name></connection>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-16.5,107,-6</points>
<intersection>-16.5 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-6,111,-6</points>
<connection>
<GID>196</GID>
<name>IN_7</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-16.5,107,-16.5</points>
<connection>
<GID>197</GID>
<name>OUT_3</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-15.5,107,-7</points>
<intersection>-15.5 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-7,111,-7</points>
<connection>
<GID>196</GID>
<name>IN_6</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-15.5,107,-15.5</points>
<connection>
<GID>197</GID>
<name>OUT_2</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 9></circuit>