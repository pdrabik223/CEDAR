<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-18.2,11.9,159.6,-80.8</PageViewport>
<gate>
<ID>2</ID>
<type>DD_KEYPAD_HEX</type>
<position>5,-12.5</position>
<output>
<ID>OUT_0</ID>161 </output>
<output>
<ID>OUT_1</ID>160 </output>
<output>
<ID>OUT_2</ID>159 </output>
<output>
<ID>OUT_3</ID>158 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>4</ID>
<type>DD_KEYPAD_HEX</type>
<position>5,-25</position>
<output>
<ID>OUT_0</ID>165 </output>
<output>
<ID>OUT_1</ID>164 </output>
<output>
<ID>OUT_2</ID>163 </output>
<output>
<ID>OUT_3</ID>162 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>6,-4</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>5,-33.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>104,-71.5</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>153 </input>
<input>
<ID>IN_3</ID>152 </input>
<input>
<ID>IN_4</ID>151 </input>
<input>
<ID>IN_5</ID>150 </input>
<input>
<ID>IN_6</ID>149 </input>
<input>
<ID>IN_7</ID>148 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 225</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>59</ID>
<type>AE_REGISTER8</type>
<position>49,-55.5</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>153 </input>
<input>
<ID>IN_3</ID>152 </input>
<input>
<ID>IN_4</ID>151 </input>
<input>
<ID>IN_5</ID>150 </input>
<input>
<ID>IN_6</ID>149 </input>
<input>
<ID>IN_7</ID>148 </input>
<output>
<ID>OUT_0</ID>144 </output>
<output>
<ID>OUT_1</ID>143 </output>
<output>
<ID>OUT_2</ID>142 </output>
<output>
<ID>OUT_3</ID>141 </output>
<output>
<ID>OUT_4</ID>140 </output>
<output>
<ID>OUT_5</ID>139 </output>
<output>
<ID>OUT_6</ID>138 </output>
<output>
<ID>OUT_7</ID>137 </output>
<input>
<ID>clear</ID>157 </input>
<input>
<ID>clock</ID>113 </input>
<input>
<ID>load</ID>145 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 225</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>61</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>26,-7</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>159 </input>
<input>
<ID>IN_2</ID>160 </input>
<input>
<ID>IN_3</ID>161 </input>
<output>
<ID>carry_out</ID>124 </output>
<input>
<ID>clear</ID>157 </input>
<input>
<ID>clock</ID>113 </input>
<input>
<ID>load</ID>108 </input>
<input>
<ID>shift_enable</ID>112 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>62</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>25.5,-24</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>164 </input>
<input>
<ID>IN_2</ID>163 </input>
<input>
<ID>IN_3</ID>162 </input>
<output>
<ID>OUT_0</ID>122 </output>
<output>
<ID>OUT_1</ID>121 </output>
<output>
<ID>OUT_2</ID>120 </output>
<output>
<ID>OUT_3</ID>119 </output>
<output>
<ID>carry_out</ID>114 </output>
<input>
<ID>clear</ID>157 </input>
<input>
<ID>clock</ID>113 </input>
<input>
<ID>load</ID>108 </input>
<input>
<ID>shift_enable</ID>111 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>63</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>25,-40</position>
<output>
<ID>OUT_0</ID>118 </output>
<output>
<ID>OUT_1</ID>117 </output>
<output>
<ID>OUT_2</ID>116 </output>
<output>
<ID>OUT_3</ID>115 </output>
<input>
<ID>carry_in</ID>114 </input>
<input>
<ID>clear</ID>157 </input>
<input>
<ID>clock</ID>113 </input>
<input>
<ID>load</ID>108 </input>
<input>
<ID>shift_enable</ID>109 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 15</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_TOGGLE</type>
<position>33,-54</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>67</ID>
<type>CC_PULSE</type>
<position>36,-54</position>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>69</ID>
<type>AE_SMALL_INVERTER</type>
<position>25,-33</position>
<input>
<ID>IN_0</ID>108 </input>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>70</ID>
<type>AE_SMALL_INVERTER</type>
<position>25.5,-17</position>
<input>
<ID>IN_0</ID>108 </input>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_SMALL_INVERTER</type>
<position>26,0</position>
<input>
<ID>IN_0</ID>108 </input>
<output>
<ID>OUT_0</ID>112 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND2</type>
<position>45,-3.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_AND2</type>
<position>46,-15</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_AND2</type>
<position>46,-20</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>120 </input>
<output>
<ID>OUT</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_AND2</type>
<position>46,-24.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_AND2</type>
<position>46,-34</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>118 </input>
<output>
<ID>OUT</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_AND2</type>
<position>46,-38</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_AND2</type>
<position>46,-42</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>116 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_AND2</type>
<position>46,-46</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_FULLADDER_4BIT</type>
<position>64.5,-8.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>143 </input>
<input>
<ID>IN_2</ID>142 </input>
<input>
<ID>IN_3</ID>141 </input>
<input>
<ID>IN_B_0</ID>125 </input>
<input>
<ID>IN_B_1</ID>126 </input>
<input>
<ID>IN_B_2</ID>127 </input>
<input>
<ID>IN_B_3</ID>128 </input>
<output>
<ID>OUT_0</ID>155 </output>
<output>
<ID>OUT_1</ID>154 </output>
<output>
<ID>OUT_2</ID>153 </output>
<output>
<ID>OUT_3</ID>152 </output>
<output>
<ID>carry_out</ID>156 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>85</ID>
<type>AE_FULLADDER_4BIT</type>
<position>64.5,-30.5</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>139 </input>
<input>
<ID>IN_2</ID>138 </input>
<input>
<ID>IN_3</ID>137 </input>
<input>
<ID>IN_B_0</ID>129 </input>
<input>
<ID>IN_B_1</ID>130 </input>
<input>
<ID>IN_B_2</ID>131 </input>
<input>
<ID>IN_B_3</ID>132 </input>
<output>
<ID>OUT_0</ID>151 </output>
<output>
<ID>OUT_1</ID>150 </output>
<output>
<ID>OUT_2</ID>149 </output>
<output>
<ID>OUT_3</ID>148 </output>
<input>
<ID>carry_in</ID>156 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>87</ID>
<type>EE_VDD</type>
<position>48.5,-47.5</position>
<output>
<ID>OUT_0</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_TOGGLE</type>
<position>33,-65.5</position>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-52,33,-1</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>-31 9</intersection>
<intersection>-17.5 4</intersection>
<intersection>-1 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>25.5,-17.5,33,-17.5</points>
<intersection>25.5 12</intersection>
<intersection>26.5 7</intersection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>26,-1,33,-1</points>
<intersection>26 13</intersection>
<intersection>27 8</intersection>
<intersection>33 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>26.5,-19,26.5,-17.5</points>
<connection>
<GID>62</GID>
<name>load</name></connection>
<intersection>-17.5 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>27,-2,27,-1</points>
<connection>
<GID>61</GID>
<name>load</name></connection>
<intersection>-1 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>25,-31,33,-31</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>26 11</intersection>
<intersection>33 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>26,-35,26,-31</points>
<connection>
<GID>63</GID>
<name>load</name></connection>
<intersection>-31 9</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>25.5,-17.5,25.5,-15</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-17.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>26,-1,26,2</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>-1 6</intersection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>25,-35,25,-35</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<connection>
<GID>63</GID>
<name>shift_enable</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-19,25.5,-19</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<connection>
<GID>62</GID>
<name>shift_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-2,26,-2</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<connection>
<GID>61</GID>
<name>shift_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-60.5,38.5,-12</points>
<intersection>-60.5 8</intersection>
<intersection>-52 9</intersection>
<intersection>-46.5 4</intersection>
<intersection>-29 3</intersection>
<intersection>-12 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-29,38.5,-29</points>
<connection>
<GID>62</GID>
<name>clock</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>26,-46.5,38.5,-46.5</points>
<intersection>26 7</intersection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>27,-12,38.5,-12</points>
<connection>
<GID>61</GID>
<name>clock</name></connection>
<intersection>38.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>26,-46.5,26,-45</points>
<connection>
<GID>63</GID>
<name>clock</name></connection>
<intersection>-46.5 4</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>38.5,-60.5,48,-60.5</points>
<connection>
<GID>59</GID>
<name>clock</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>36,-52,38.5,-52</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-35,22.5,-29</points>
<intersection>-35 4</intersection>
<intersection>-29 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>22.5,-29,24,-29</points>
<connection>
<GID>62</GID>
<name>carry_out</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>22.5,-35,23.5,-35</points>
<connection>
<GID>63</GID>
<name>carry_in</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-47,34,-41.5</points>
<intersection>-47 2</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-41.5,34,-41.5</points>
<connection>
<GID>63</GID>
<name>OUT_3</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-47,43,-47</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-43,35.5,-40.5</points>
<intersection>-43 2</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-40.5,35.5,-40.5</points>
<connection>
<GID>63</GID>
<name>OUT_2</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-43,43,-43</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-39.5,35.5,-39</points>
<intersection>-39.5 1</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-39.5,35.5,-39.5</points>
<connection>
<GID>63</GID>
<name>OUT_1</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-39,43,-39</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-38.5,35.5,-35</points>
<intersection>-38.5 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-38.5,35.5,-38.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-35,43,-35</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-25.5,43,-25.5</points>
<connection>
<GID>62</GID>
<name>OUT_3</name></connection>
<connection>
<GID>76</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-24.5,36,-21</points>
<intersection>-24.5 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-24.5,36,-24.5</points>
<connection>
<GID>62</GID>
<name>OUT_2</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-21,43,-21</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-23.5,34.5,-16</points>
<intersection>-23.5 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-23.5,34.5,-23.5</points>
<connection>
<GID>62</GID>
<name>OUT_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-16,43,-16</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-22.5,35,-4.5</points>
<intersection>-22.5 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-22.5,35,-22.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-4.5,42,-4.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-14,24.5,-12</points>
<connection>
<GID>61</GID>
<name>carry_out</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-14,43,-14</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection>
<intersection>40 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>40,-45,40,-2.5</points>
<intersection>-45 26</intersection>
<intersection>-41 31</intersection>
<intersection>-37 30</intersection>
<intersection>-33 29</intersection>
<intersection>-23.5 3</intersection>
<intersection>-19 6</intersection>
<intersection>-14 1</intersection>
<intersection>-2.5 28</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>40,-23.5,43,-23.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>40 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>40,-19,43,-19</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>40 2</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>40,-45,43,-45</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>40 2</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>40,-2.5,42,-2.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>40 2</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>40,-33,43,-33</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>40 2</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>40,-37,43,-37</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>40 2</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>40,-41,43,-41</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>40 2</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3.5,60.5,-3.5</points>
<connection>
<GID>84</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>73</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-15,52.5,-4.5</points>
<intersection>-15 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-4.5,60.5,-4.5</points>
<connection>
<GID>84</GID>
<name>IN_B_1</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-15,52.5,-15</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-20,53.5,-5.5</points>
<intersection>-20 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-20,53.5,-20</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-5.5,60.5,-5.5</points>
<connection>
<GID>84</GID>
<name>IN_B_2</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-24.5,54.5,-6.5</points>
<intersection>-24.5 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-6.5,60.5,-6.5</points>
<connection>
<GID>84</GID>
<name>IN_B_3</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-24.5,54.5,-24.5</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-34,52,-25.5</points>
<intersection>-34 1</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-34,52,-34</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-25.5,60.5,-25.5</points>
<connection>
<GID>85</GID>
<name>IN_B_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-38,51,-26.5</points>
<intersection>-38 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-38,51,-38</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-26.5,60.5,-26.5</points>
<connection>
<GID>85</GID>
<name>IN_B_1</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-42,53,-27.5</points>
<intersection>-42 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-42,53,-42</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-27.5,60.5,-27.5</points>
<connection>
<GID>85</GID>
<name>IN_B_2</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-46,54,-28.5</points>
<intersection>-46 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-46,54,-46</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-28.5,60.5,-28.5</points>
<connection>
<GID>85</GID>
<name>IN_B_3</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-48.5,60.5,-48.5</points>
<intersection>53 3</intersection>
<intersection>60.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>53,-51.5,53,-48.5</points>
<connection>
<GID>59</GID>
<name>OUT_7</name></connection>
<intersection>-48.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>60.5,-48.5,60.5,-35.5</points>
<connection>
<GID>85</GID>
<name>IN_3</name></connection>
<intersection>-48.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-52.5,56.5,-34.5</points>
<intersection>-52.5 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-52.5,56.5,-52.5</points>
<connection>
<GID>59</GID>
<name>OUT_6</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-34.5,60.5,-34.5</points>
<connection>
<GID>85</GID>
<name>IN_2</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-53.5,57,-33.5</points>
<intersection>-53.5 1</intersection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-53.5,57,-53.5</points>
<connection>
<GID>59</GID>
<name>OUT_5</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-33.5,60.5,-33.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-54.5,55.5,-32.5</points>
<intersection>-54.5 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-54.5,55.5,-54.5</points>
<connection>
<GID>59</GID>
<name>OUT_4</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-32.5,60.5,-32.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-55.5,59.5,-13.5</points>
<intersection>-55.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-55.5,59.5,-55.5</points>
<connection>
<GID>59</GID>
<name>OUT_3</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59.5,-13.5,60.5,-13.5</points>
<connection>
<GID>84</GID>
<name>IN_3</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-56.5,58.5,-12.5</points>
<intersection>-56.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-56.5,58.5,-56.5</points>
<connection>
<GID>59</GID>
<name>OUT_2</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58.5,-12.5,60.5,-12.5</points>
<connection>
<GID>84</GID>
<name>IN_2</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-57.5,57.5,-11.5</points>
<intersection>-57.5 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-57.5,57.5,-57.5</points>
<connection>
<GID>59</GID>
<name>OUT_1</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-11.5,60.5,-11.5</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-58.5,56,-10.5</points>
<intersection>-58.5 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-58.5,56,-58.5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-10.5,60.5,-10.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-49.5,48,-48.5</points>
<connection>
<GID>59</GID>
<name>load</name></connection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-48.5,48.5,-48.5</points>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>82,-67.5,82,-32</points>
<intersection>-67.5 5</intersection>
<intersection>-32 13</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>39.5,-67.5,99,-67.5</points>
<connection>
<GID>57</GID>
<name>IN_7</name></connection>
<intersection>39.5 8</intersection>
<intersection>82 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>39.5,-67.5,39.5,-51.5</points>
<intersection>-67.5 5</intersection>
<intersection>-51.5 14</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>68.5,-32,82,-32</points>
<connection>
<GID>85</GID>
<name>OUT_3</name></connection>
<intersection>82 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>39.5,-51.5,45,-51.5</points>
<connection>
<GID>59</GID>
<name>IN_7</name></connection>
<intersection>39.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-68.5,79.5,-31</points>
<intersection>-68.5 1</intersection>
<intersection>-31 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-68.5,99,-68.5</points>
<connection>
<GID>57</GID>
<name>IN_6</name></connection>
<intersection>42.5 6</intersection>
<intersection>79.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>42.5,-68.5,42.5,-52.5</points>
<intersection>-68.5 1</intersection>
<intersection>-52.5 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-31,79.5,-31</points>
<connection>
<GID>85</GID>
<name>OUT_2</name></connection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>42.5,-52.5,45,-52.5</points>
<connection>
<GID>59</GID>
<name>IN_6</name></connection>
<intersection>42.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-69.5,76.5,-30</points>
<intersection>-69.5 1</intersection>
<intersection>-30 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-69.5,99,-69.5</points>
<connection>
<GID>57</GID>
<name>IN_5</name></connection>
<intersection>41.5 6</intersection>
<intersection>76.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>41.5,-69.5,41.5,-53.5</points>
<intersection>-69.5 1</intersection>
<intersection>-53.5 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-30,76.5,-30</points>
<connection>
<GID>85</GID>
<name>OUT_1</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>41.5,-53.5,45,-53.5</points>
<connection>
<GID>59</GID>
<name>IN_5</name></connection>
<intersection>41.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-70.5,73.5,-29</points>
<intersection>-70.5 1</intersection>
<intersection>-29 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-70.5,99,-70.5</points>
<connection>
<GID>57</GID>
<name>IN_4</name></connection>
<intersection>44 6</intersection>
<intersection>73.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>44,-70.5,44,-54.5</points>
<intersection>-70.5 1</intersection>
<intersection>-54.5 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-29,73.5,-29</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>44,-54.5,45,-54.5</points>
<connection>
<GID>59</GID>
<name>IN_4</name></connection>
<intersection>44 6</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-71.5,87.5,-10</points>
<intersection>-71.5 1</intersection>
<intersection>-10 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-71.5,99,-71.5</points>
<connection>
<GID>57</GID>
<name>IN_3</name></connection>
<intersection>44.5 6</intersection>
<intersection>87.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>44.5,-71.5,44.5,-55.5</points>
<intersection>-71.5 1</intersection>
<intersection>-55.5 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-10,87.5,-10</points>
<connection>
<GID>84</GID>
<name>OUT_3</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>44.5,-55.5,45,-55.5</points>
<connection>
<GID>59</GID>
<name>IN_3</name></connection>
<intersection>44.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-72.5,89,-9</points>
<intersection>-72.5 1</intersection>
<intersection>-9 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-72.5,99,-72.5</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<intersection>45 6</intersection>
<intersection>89 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>45,-72.5,45,-56.5</points>
<connection>
<GID>59</GID>
<name>IN_2</name></connection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-9,89,-9</points>
<connection>
<GID>84</GID>
<name>OUT_2</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-73.5,90.5,-8</points>
<intersection>-73.5 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-73.5,99,-73.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>43 8</intersection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-8,90.5,-8</points>
<connection>
<GID>84</GID>
<name>OUT_1</name></connection>
<intersection>90.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>43,-73.5,43,-57.5</points>
<intersection>-73.5 1</intersection>
<intersection>-57.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>43,-57.5,45,-57.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>43 8</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-74.5,92,-7</points>
<intersection>-74.5 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-74.5,99,-74.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>40.5 7</intersection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-7,92,-7</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>92 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>40.5,-74.5,40.5,-58.5</points>
<intersection>-74.5 1</intersection>
<intersection>-58.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>40.5,-58.5,45,-58.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>40.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-22.5,63.5,-16.5</points>
<connection>
<GID>84</GID>
<name>carry_out</name></connection>
<connection>
<GID>85</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-63.5,33,-58.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<intersection>-62 2</intersection>
<intersection>-58.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50,-62,50,-60.5</points>
<connection>
<GID>59</GID>
<name>clear</name></connection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>33,-62,50,-62</points>
<intersection>33 0</intersection>
<intersection>50 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-58.5,33,-58.5</points>
<intersection>30.5 4</intersection>
<intersection>33 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-58.5,30.5,-29</points>
<intersection>-58.5 3</intersection>
<intersection>-45 6</intersection>
<intersection>-29 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>25.5,-29,31,-29</points>
<connection>
<GID>62</GID>
<name>clear</name></connection>
<intersection>30.5 4</intersection>
<intersection>31 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>25,-45,30.5,-45</points>
<connection>
<GID>63</GID>
<name>clear</name></connection>
<intersection>30.5 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>31,-29,31,-12</points>
<intersection>-29 5</intersection>
<intersection>-12 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>26,-12,31,-12</points>
<connection>
<GID>61</GID>
<name>clear</name></connection>
<intersection>31 7</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-9.5,16,-5.5</points>
<intersection>-9.5 2</intersection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-5.5,22.5,-5.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-9.5,16,-9.5</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-11.5,16,-6.5</points>
<intersection>-11.5 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-6.5,22.5,-6.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-11.5,16,-11.5</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-13.5,16,-7.5</points>
<intersection>-13.5 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-13.5,16,-13.5</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-7.5,22.5,-7.5</points>
<connection>
<GID>61</GID>
<name>IN_2</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-15.5,16,-8.5</points>
<intersection>-15.5 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-15.5,16,-15.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-8.5,22.5,-8.5</points>
<connection>
<GID>61</GID>
<name>IN_3</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-25.5,16,-22</points>
<intersection>-25.5 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-25.5,22,-25.5</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-22,16,-22</points>
<connection>
<GID>4</GID>
<name>OUT_3</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-24.5,16,-24</points>
<intersection>-24.5 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-24.5,22,-24.5</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-24,16,-24</points>
<connection>
<GID>4</GID>
<name>OUT_2</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-26,16,-23.5</points>
<intersection>-26 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-23.5,22,-23.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-26,16,-26</points>
<connection>
<GID>4</GID>
<name>OUT_1</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-28,16,-22.5</points>
<intersection>-28 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-22.5,22,-22.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-28,16,-28</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 9></circuit>