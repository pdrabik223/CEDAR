<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-49.1106,-62.2952,55.3551,-179.819</PageViewport>
<gate>
<ID>2</ID>
<type>BA_NAND2</type>
<position>1.5,15.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>0,22</position>
<gparam>LABEL_TEXT tabela 5-1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>0,1.5</position>
<gparam>LABEL_TEXT tabela 5-2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>-1,-20</position>
<gparam>LABEL_TEXT tabela 5-3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>-6.5,16.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>-3.5,-41.5</position>
<gparam>LABEL_TEXT tabela 5-4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>-8.5,-55.5</position>
<gparam>LABEL_TEXT sumator niezupe�ny</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>-4,-73</position>
<gparam>LABEL_TEXT niezupe�ny uk�ad r�nicy</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>-13.5,16.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>-8.5,-97</position>
<gparam>LABEL_TEXT Uk�ad por�wnuj�cy binarnie</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>-14,8.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_SMALL_INVERTER</type>
<position>6.5,15.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_SMALL_INVERTER</type>
<position>6.5,9.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>15</ID>
<type>BA_NAND2</type>
<position>1.5,9.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_SMALL_INVERTER</type>
<position>-6,8.5</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>-7,-139</position>
<gparam>LABEL_TEXT Uk�ad kontroli parzysto�ci</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>BE_NOR2</type>
<position>13,13</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_SMALL_INVERTER</type>
<position>26,13</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>29,13</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>BE_NOR2</type>
<position>2,-4.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>BE_NOR2</type>
<position>1.5,-11</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>BE_NOR2</type>
<position>17,-8.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_SMALL_INVERTER</type>
<position>-3.5,-10</position>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_SMALL_INVERTER</type>
<position>-3.5,-12</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>23,-8.5</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>-13.5,-8.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>-13.5,-3.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>BA_NAND2</type>
<position>-2.5,-31</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_SMALL_INVERTER</type>
<position>2.5,-31</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>32</ID>
<type>BE_NOR2</type>
<position>7.5,-30</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>12,-30</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>BE_NOR2</type>
<position>1,-25.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>-13.5,-32</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>-13.5,-24.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>-13.5,-49</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>-13.5,-47</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>-16,-144</position>
<gparam>LABEL_TEXT B4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AI_XOR2</type>
<position>-5.5,-48</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>GA_LED</type>
<position>14.5,-48</position>
<input>
<ID>N_in0</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>-16,-146.5</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>-16,-150.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>BA_NAND2</type>
<position>-7.5,-67.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_SMALL_INVERTER</type>
<position>-2.5,-67.5</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>7.5,-62</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>7.5,-67.5</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>-19,-68.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>-19,-61</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AI_XOR2</type>
<position>-7,-62</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>-16,-155</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>BA_NAND2</type>
<position>-7.5,-84</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>-16,-160</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>7.5,-79</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>GA_LED</type>
<position>9.5,-87</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>-20,-86</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>-20,-78</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>58</ID>
<type>AI_XOR2</type>
<position>-7,-79</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>BA_NAND2</type>
<position>-1.5,-85.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>BA_NAND2</type>
<position>4.5,-87</position>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>AI_XOR2</type>
<position>-7,-110</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_SMALL_INVERTER</type>
<position>-2,-110</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>2.5,-159</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AI_XOR2</type>
<position>-7,-115.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>AE_SMALL_INVERTER</type>
<position>-2,-115.5</position>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AI_XOR2</type>
<position>-7,-121</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>AE_SMALL_INVERTER</type>
<position>-2,-121</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>68</ID>
<type>AI_XOR2</type>
<position>-7,-126.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_SMALL_INVERTER</type>
<position>-2,-126.5</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>-17.5,17</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_AND4</type>
<position>9.5,-118.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>51 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>-20,-104</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>-17.5,-104</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>-15,-104</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>-12.5,-104</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>-17.5,9</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>31.5,13.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>-16.5,-3</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>-16.5,-8</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>-19.5,-130.5</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_TOGGLE</type>
<position>-17,-130.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>-14.5,-130.5</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_TOGGLE</type>
<position>-12,-130.5</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>13.5,-118.5</position>
<input>
<ID>N_in0</ID>61 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_TOGGLE</type>
<position>-12.5,-144.5</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>-12.5,-146.5</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_TOGGLE</type>
<position>-12.5,-151</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_TOGGLE</type>
<position>-12.5,-155.5</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_TOGGLE</type>
<position>-12.5,-160.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>90</ID>
<type>AI_XOR2</type>
<position>-4.5,-145.5</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AI_XOR2</type>
<position>-4.5,-150</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AI_XOR2</type>
<position>-4.5,-154.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AI_XOR2</type>
<position>-4.5,-159.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>-0.5,-159.5</position>
<input>
<ID>N_in0</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>25,-8</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>-17,-24</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>-16.5,-31.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>14.5,-29.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>17,-47.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>-17,-46.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>-17,-49</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>-22.5,-60.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>-22.5,-68</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>10.5,-61</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>10.5,-67</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>-23,-77.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>-23,-85</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>13,-79</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>13,-86.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>-22.5,-100.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>-18.5,-100.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>-14.5,-100.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>-10.5,-100.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>-22.5,-133</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>-18.5,-133</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>-14.5,-133</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>-10.5,-133</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>22.5,-118</position>
<gparam>LABEL_TEXT true/false</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>GA_LED</type>
<position>19.5,13</position>
<input>
<ID>N_in0</ID>4 </input>
<input>
<ID>N_in1</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>19.5,16</position>
<gparam>LABEL_TEXT !X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4.5,16.5,-1.5,16.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,13,24,13</points>
<connection>
<GID>119</GID>
<name>N_in1</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-11.5,16.5,-8.5,16.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-10 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-10,10.5,-10,16.5</points>
<intersection>10.5 3</intersection>
<intersection>16.5 0</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-10,10.5,-1.5,10.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-10 2</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,13,18.5,13</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>119</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,15.5,4.5,15.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>13</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,9.5,4.5,9.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>15</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4,8.5,-1.5,8.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,8.5,-8,8.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-9 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-9,8.5,-9,14.5</points>
<intersection>8.5 1</intersection>
<intersection>14.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-9,14.5,-1.5,14.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-9 3</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,14,9,15.5</points>
<intersection>14 2</intersection>
<intersection>15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,15.5,9,15.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9,14,10,14</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,9.5,9,12</points>
<intersection>9.5 1</intersection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,9.5,9,9.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9,12,10,12</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,13,28,13</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<connection>
<GID>21</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-10,-1.5,-10</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-12,-1.5,-12</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-11,9,-9.5</points>
<intersection>-11 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-9.5,14,-9.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-11,9,-11</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-7.5,9.5,-4.5</points>
<intersection>-7.5 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-4.5,9.5,-4.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-7.5,14,-7.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-8.5,22,-8.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<connection>
<GID>27</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-10,-8,-3.5</points>
<intersection>-10 5</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11.5,-3.5,-1,-3.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>-8 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-8,-10,-5.5,-10</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-12,-10,-5.5</points>
<intersection>-12 3</intersection>
<intersection>-8.5 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11.5,-8.5,-10,-8.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10,-5.5,-1,-5.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-10,-12,-5.5,-12</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-31,0.5,-31</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<connection>
<GID>31</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-31,4.5,-31</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>10.5,-30,11,-30</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<connection>
<GID>33</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-29,4,-25.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-29,4.5,-29</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-32,-5.5,-32</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>-10 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-10,-32,-10,-26.5</points>
<intersection>-32 1</intersection>
<intersection>-26.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-10,-26.5,-2,-26.5</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>-10 4</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9,-30,-9,-24.5</points>
<intersection>-30 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9,-30,-5.5,-30</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11.5,-24.5,-2,-24.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>-9 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-49,-8.5,-49</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-47,-8.5,-47</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2.5,-48,13.5,-48</points>
<connection>
<GID>41</GID>
<name>N_in0</name></connection>
<connection>
<GID>40</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-4.5,-67.5,-4.5,-67.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-67.5,6.5,-67.5</points>
<connection>
<GID>47</GID>
<name>N_in0</name></connection>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17,-68.5,-10.5,-68.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-12 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-12,-68.5,-12,-63</points>
<intersection>-68.5 1</intersection>
<intersection>-63 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-12,-63,-10,-63</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-12 8</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-66.5,-13.5,-61</points>
<intersection>-66.5 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,-61,-10,-61</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,-66.5,-10.5,-66.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4,-62,6.5,-62</points>
<connection>
<GID>46</GID>
<name>N_in0</name></connection>
<connection>
<GID>50</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-83,-13.5,-78</points>
<intersection>-83 2</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-18,-78,-10,-78</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,-83,-10.5,-83</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4,-79,6.5,-79</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<connection>
<GID>54</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-84.5,-4.5,-84</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-86,1.5,-85.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<connection>
<GID>59</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>7.5,-87,8.5,-87</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<connection>
<GID>55</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18,-86,-4.5,-86</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>-12 4</intersection>
<intersection>-4.5 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12,-86,-12,-80</points>
<intersection>-86 1</intersection>
<intersection>-80 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-12,-80,-10,-80</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>-12 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-4.5,-86.5,-4.5,-86</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>-86 1</intersection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-110,-4,-110</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<connection>
<GID>62</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-115.5,-4,-115.5</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<connection>
<GID>65</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-121,-4,-121</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-126.5,-4,-126.5</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<connection>
<GID>69</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-115.5,5,-110</points>
<intersection>-115.5 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-110,5,-110</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-115.5,6.5,-115.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-117.5,3,-115.5</points>
<intersection>-117.5 2</intersection>
<intersection>-115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-115.5,3,-115.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-117.5,6.5,-117.5</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-121,3,-119.5</points>
<intersection>-121 1</intersection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-121,3,-121</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-119.5,6.5,-119.5</points>
<connection>
<GID>71</GID>
<name>IN_2</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-126.5,5,-121.5</points>
<intersection>-126.5 1</intersection>
<intersection>-121.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-126.5,5,-126.5</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-121.5,6.5,-121.5</points>
<connection>
<GID>71</GID>
<name>IN_3</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-128.5,-12,-127.5</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,-127.5,-10,-127.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,-125.5,-20,-106</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20,-125.5,-10,-125.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>-20 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-128.5,-14.5,-122</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>-122 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-122,-10,-122</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-120,-10,-120</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-17.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-17.5,-120,-17.5,-106</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>-120 1</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-128.5,-16,-116.5</points>
<intersection>-128.5 2</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-116.5,-10,-116.5</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-17,-128.5,-16,-128.5</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,-114.5,-15,-106</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>-114.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-114.5,-10,-114.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19,-128.5,-19,-111</points>
<intersection>-128.5 2</intersection>
<intersection>-111 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19,-111,-10,-111</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>-19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-128.5,-19,-128.5</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>-19 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-109,-12.5,-106</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,-109,-10,-109</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-118.5,12.5,-118.5</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<connection>
<GID>84</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-157,1.5,-154.5</points>
<intersection>-157 1</intersection>
<intersection>-154.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-157,1.5,-157</points>
<intersection>-7.5 3</intersection>
<intersection>1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,-154.5,1.5,-154.5</points>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>1.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-7.5,-158.5,-7.5,-157</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>-157 1</intersection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-152,2,-150</points>
<intersection>-152 2</intersection>
<intersection>-150 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,-150,2,-150</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-152,2,-152</points>
<intersection>-7.5 3</intersection>
<intersection>2 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-7.5,-153.5,-7.5,-152</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>-152 2</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-148,2,-145.5</points>
<intersection>-148 2</intersection>
<intersection>-145.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,-145.5,2,-145.5</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-148,2,-148</points>
<intersection>-7.5 3</intersection>
<intersection>2 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-7.5,-149,-7.5,-148</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-148 2</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-146.5,-7.5,-146.5</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<connection>
<GID>90</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-144.5,-7.5,-144.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-151,-7.5,-151</points>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<connection>
<GID>91</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-155.5,-7.5,-155.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<connection>
<GID>92</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-160.5,-7.5,-160.5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-7.5,-160.5,-7.5,-160.5</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>-160.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-159.5,-1.5,-159.5</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<connection>
<GID>94</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-2.11928e-006,0,81.6,-91.8</PageViewport></page 1>
<page 2>
<PageViewport>-2.11928e-006,0,81.6,-91.8</PageViewport></page 2>
<page 3>
<PageViewport>-2.11928e-006,0,81.6,-91.8</PageViewport></page 3>
<page 4>
<PageViewport>-2.11928e-006,0,81.6,-91.8</PageViewport></page 4>
<page 5>
<PageViewport>-2.11928e-006,0,81.6,-91.8</PageViewport></page 5>
<page 6>
<PageViewport>-2.11928e-006,0,81.6,-91.8</PageViewport></page 6>
<page 7>
<PageViewport>-2.11928e-006,0,81.6,-91.8</PageViewport></page 7>
<page 8>
<PageViewport>-2.11928e-006,0,81.6,-91.8</PageViewport></page 8>
<page 9>
<PageViewport>-2.11928e-006,0,81.6,-91.8</PageViewport></page 9></circuit>