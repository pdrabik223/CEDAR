<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-153.854,50.4876,193.112,-121.011</PageViewport>
<gate>
<ID>2</ID>
<type>DD_KEYPAD_HEX</type>
<position>7,-29.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<output>
<ID>OUT_1</ID>16 </output>
<output>
<ID>OUT_2</ID>17 </output>
<output>
<ID>OUT_3</ID>18 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 13</lparam></gate>
<gate>
<ID>4</ID>
<type>GA_LED</type>
<position>4.5,-48</position>
<input>
<ID>N_in1</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>GA_LED</type>
<position>6.5,-48</position>
<input>
<ID>N_in0</ID>1 </input>
<input>
<ID>N_in1</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>8.5,-48</position>
<input>
<ID>N_in0</ID>2 </input>
<input>
<ID>N_in1</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>4.5,-40</position>
<input>
<ID>N_in1</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>6.5,-40</position>
<input>
<ID>N_in0</ID>3 </input>
<input>
<ID>N_in1</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>8.5,-40</position>
<input>
<ID>N_in0</ID>4 </input>
<input>
<ID>N_in1</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>4.5,-56</position>
<input>
<ID>N_in1</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>6.5,-56</position>
<input>
<ID>N_in0</ID>5 </input>
<input>
<ID>N_in1</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>8.5,-56</position>
<input>
<ID>N_in0</ID>6 </input>
<input>
<ID>N_in1</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>GA_LED</type>
<position>10.5,-42</position>
<input>
<ID>N_in1</ID>43 </input>
<input>
<ID>N_in2</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>10.5,-44</position>
<input>
<ID>N_in2</ID>8 </input>
<input>
<ID>N_in3</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>GA_LED</type>
<position>10.5,-46</position>
<input>
<ID>N_in3</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>2.5,-42</position>
<input>
<ID>N_in2</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>2.5,-44</position>
<input>
<ID>N_in1</ID>47 </input>
<input>
<ID>N_in2</ID>10 </input>
<input>
<ID>N_in3</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>2.5,-46</position>
<input>
<ID>N_in3</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>10.5,-50</position>
<input>
<ID>N_in1</ID>44 </input>
<input>
<ID>N_in2</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>10.5,-52</position>
<input>
<ID>N_in2</ID>12 </input>
<input>
<ID>N_in3</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>10.5,-54</position>
<input>
<ID>N_in3</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>GA_LED</type>
<position>2.5,-50</position>
<input>
<ID>N_in2</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>2.5,-52</position>
<input>
<ID>N_in1</ID>46 </input>
<input>
<ID>N_in2</ID>14 </input>
<input>
<ID>N_in3</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>2.5,-54</position>
<input>
<ID>N_in3</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>BE_ROM_8x8</type>
<position>27.5,-29</position>
<input>
<ID>ADDRESS_0</ID>19 </input>
<input>
<ID>ADDRESS_1</ID>31 </input>
<input>
<ID>ADDRESS_2</ID>32 </input>
<input>
<ID>ADDRESS_3</ID>34 </input>
<output>
<ID>DATA_OUT_0</ID>35 </output>
<output>
<ID>DATA_OUT_1</ID>36 </output>
<output>
<ID>DATA_OUT_2</ID>37 </output>
<output>
<ID>DATA_OUT_3</ID>38 </output>
<output>
<ID>DATA_OUT_4</ID>39 </output>
<output>
<ID>DATA_OUT_5</ID>40 </output>
<output>
<ID>DATA_OUT_6</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:0 63</lparam>
<lparam>Address:1 6</lparam>
<lparam>Address:2 91</lparam>
<lparam>Address:3 79</lparam>
<lparam>Address:4 102</lparam>
<lparam>Address:5 109</lparam>
<lparam>Address:6 125</lparam>
<lparam>Address:7 7</lparam>
<lparam>Address:8 127</lparam>
<lparam>Address:9 103</lparam>
<lparam>Address:10 119</lparam>
<lparam>Address:11 124</lparam>
<lparam>Address:12 57</lparam>
<lparam>Address:13 94</lparam>
<lparam>Address:14 121</lparam>
<lparam>Address:15 113</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>13,-32.5</position>
<input>
<ID>N_in0</ID>15 </input>
<input>
<ID>N_in1</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>15,-30.5</position>
<input>
<ID>N_in0</ID>16 </input>
<input>
<ID>N_in1</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>17,-28.5</position>
<input>
<ID>N_in0</ID>17 </input>
<input>
<ID>N_in1</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>19,-26.5</position>
<input>
<ID>N_in0</ID>18 </input>
<input>
<ID>N_in1</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>GA_LED</type>
<position>32,-40</position>
<input>
<ID>N_in0</ID>42 </input>
<input>
<ID>N_in3</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>30,-42</position>
<input>
<ID>N_in0</ID>43 </input>
<input>
<ID>N_in3</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>28,-44</position>
<input>
<ID>N_in0</ID>44 </input>
<input>
<ID>N_in3</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>GA_LED</type>
<position>26,-46</position>
<input>
<ID>N_in0</ID>45 </input>
<input>
<ID>N_in3</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>24,-48</position>
<input>
<ID>N_in0</ID>46 </input>
<input>
<ID>N_in3</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>GA_LED</type>
<position>22,-50</position>
<input>
<ID>N_in0</ID>47 </input>
<input>
<ID>N_in3</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>20,-52</position>
<input>
<ID>N_in0</ID>48 </input>
<input>
<ID>N_in3</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>6.5,-36.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>13,-43.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>13,-51</position>
<gparam>LABEL_TEXT c</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>6.5,-58</position>
<gparam>LABEL_TEXT d</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>0,-51.5</position>
<gparam>LABEL_TEXT e</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>6.5,-45.5</position>
<gparam>LABEL_TEXT g</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-48,5.5,-48</points>
<connection>
<GID>4</GID>
<name>N_in1</name></connection>
<connection>
<GID>7</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-48,7.5,-48</points>
<connection>
<GID>7</GID>
<name>N_in1</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-40,5.5,-40</points>
<connection>
<GID>9</GID>
<name>N_in1</name></connection>
<connection>
<GID>10</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-40,7.5,-40</points>
<connection>
<GID>10</GID>
<name>N_in1</name></connection>
<connection>
<GID>11</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>5.5,-56,5.5,-56</points>
<connection>
<GID>12</GID>
<name>N_in1</name></connection>
<connection>
<GID>13</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-56,7.5,-56</points>
<connection>
<GID>13</GID>
<name>N_in1</name></connection>
<connection>
<GID>14</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>10.5,-43,10.5,-43</points>
<connection>
<GID>15</GID>
<name>N_in2</name></connection>
<connection>
<GID>16</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>10.5,-45,10.5,-45</points>
<connection>
<GID>16</GID>
<name>N_in2</name></connection>
<connection>
<GID>17</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>2.5,-43,2.5,-43</points>
<connection>
<GID>19</GID>
<name>N_in2</name></connection>
<connection>
<GID>20</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>2.5,-45,2.5,-45</points>
<connection>
<GID>20</GID>
<name>N_in2</name></connection>
<connection>
<GID>21</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>10.5,-51,10.5,-51</points>
<connection>
<GID>22</GID>
<name>N_in2</name></connection>
<connection>
<GID>23</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>10.5,-53,10.5,-53</points>
<connection>
<GID>23</GID>
<name>N_in2</name></connection>
<connection>
<GID>24</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>2.5,-51,2.5,-51</points>
<connection>
<GID>25</GID>
<name>N_in2</name></connection>
<connection>
<GID>26</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>2.5,-53,2.5,-53</points>
<connection>
<GID>26</GID>
<name>N_in2</name></connection>
<connection>
<GID>27</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-32.5,12,-32.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>33</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-30.5,14,-30.5</points>
<connection>
<GID>35</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-28.5,16,-28.5</points>
<connection>
<GID>37</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-26.5,18,-26.5</points>
<connection>
<GID>39</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-32.5,22.5,-32.5</points>
<connection>
<GID>29</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>33</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-31.5,19,-30.5</points>
<intersection>-31.5 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-30.5,19,-30.5</points>
<connection>
<GID>35</GID>
<name>N_in1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-31.5,22.5,-31.5</points>
<connection>
<GID>29</GID>
<name>ADDRESS_1</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-30.5,20,-28.5</points>
<intersection>-30.5 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-30.5,22.5,-30.5</points>
<connection>
<GID>29</GID>
<name>ADDRESS_2</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-28.5,20,-28.5</points>
<connection>
<GID>37</GID>
<name>N_in1</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-29.5,21,-26.5</points>
<intersection>-29.5 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-26.5,21,-26.5</points>
<connection>
<GID>39</GID>
<name>N_in1</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-29.5,22.5,-29.5</points>
<connection>
<GID>29</GID>
<name>ADDRESS_3</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-39,32,-36</points>
<connection>
<GID>41</GID>
<name>N_in3</name></connection>
<intersection>-36 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>31,-36,32,-36</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-41,30,-36</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>59</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-43,28,-38.5</points>
<connection>
<GID>60</GID>
<name>N_in3</name></connection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>28,-38.5,29,-38.5</points>
<intersection>28 0</intersection>
<intersection>29 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>29,-38.5,29,-36</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-38.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-45,26,-38</points>
<connection>
<GID>61</GID>
<name>N_in3</name></connection>
<intersection>-38 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>28,-38,28,-36</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>26,-38,28,-38</points>
<intersection>26 0</intersection>
<intersection>28 1</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-47,24,-37.5</points>
<connection>
<GID>62</GID>
<name>N_in3</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>27,-37.5,27,-36</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_4</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24,-37.5,27,-37.5</points>
<intersection>24 0</intersection>
<intersection>27 1</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-49,22,-37</points>
<connection>
<GID>63</GID>
<name>N_in3</name></connection>
<intersection>-37 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>26,-37,26,-36</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_5</name></connection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22,-37,26,-37</points>
<intersection>22 0</intersection>
<intersection>26 1</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-51,20,-36.5</points>
<connection>
<GID>64</GID>
<name>N_in3</name></connection>
<intersection>-36.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>20,-36.5,25,-36.5</points>
<intersection>20 0</intersection>
<intersection>25 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>25,-36.5,25,-36</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_6</name></connection>
<intersection>-36.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9.5,-40,31,-40</points>
<connection>
<GID>41</GID>
<name>N_in0</name></connection>
<connection>
<GID>11</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-42,29,-42</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<connection>
<GID>15</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-50,14,-44</points>
<intersection>-50 1</intersection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-50,14,-50</points>
<connection>
<GID>22</GID>
<name>N_in1</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-44,27,-44</points>
<connection>
<GID>60</GID>
<name>N_in0</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-56,15.5,-46</points>
<intersection>-56 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-56,15.5,-56</points>
<connection>
<GID>14</GID>
<name>N_in1</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-46,25,-46</points>
<connection>
<GID>61</GID>
<name>N_in0</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-57.5,15,-48</points>
<intersection>-57.5 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-57.5,15,-57.5</points>
<intersection>3.5 3</intersection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-48,23,-48</points>
<connection>
<GID>62</GID>
<name>N_in0</name></connection>
<intersection>15 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>3.5,-57.5,3.5,-52</points>
<connection>
<GID>26</GID>
<name>N_in1</name></connection>
<intersection>-57.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-57.5,12.5,-50</points>
<intersection>-57.5 1</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-57.5,12.5,-57.5</points>
<intersection>3.5 3</intersection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-50,21,-50</points>
<connection>
<GID>63</GID>
<name>N_in0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>3.5,-57.5,3.5,-44</points>
<connection>
<GID>20</GID>
<name>N_in1</name></connection>
<intersection>-57.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-56.5,18,-52</points>
<intersection>-56.5 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-56.5,18,-56.5</points>
<intersection>9.5 3</intersection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-52,19,-52</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<intersection>18 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>9.5,-56.5,9.5,-48</points>
<connection>
<GID>8</GID>
<name>N_in1</name></connection>
<intersection>-56.5 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 1>
<page 2>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 2>
<page 3>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 3>
<page 4>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 4>
<page 5>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 5>
<page 6>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 6>
<page 7>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 7>
<page 8>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 8>
<page 9>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 9></circuit>