<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-9.01138,1.99554,53.4499,-63.1508</PageViewport></page 0>
<page 1>
<PageViewport>-37.7298,45.6002,61.4011,-57.792</PageViewport>
<gate>
<ID>1</ID>
<type>BM_NORX2</type>
<position>101,-7</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>GA_LED</type>
<position>12,-11</position>
<gparam>LED_BOX -30,-20,30,20</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AE_OR3</type>
<position>113,51.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>4</ID>
<type>GA_LED</type>
<position>1.5,-41</position>
<gparam>LED_BOX -30,-20,30,20</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AE_SMALL_INVERTER</type>
<position>108,53.5</position>
<input>
<ID>IN_0</ID>134 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>BM_NORX2</type>
<position>107,50.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>DA_FROM</type>
<position>22,-6</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>9</ID>
<type>DA_FROM</type>
<position>23.5,4</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID .</lparam></gate>
<gate>
<ID>10</ID>
<type>DA_FROM</type>
<position>32,-5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>11</ID>
<type>DA_FROM</type>
<position>23.5,-9</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID '</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND3</type>
<position>101.5,-23.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>133 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>14</ID>
<type>DA_FROM</type>
<position>22,-19</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID 2</lparam></gate>
<gate>
<ID>15</ID>
<type>DA_FROM</type>
<position>32,-19</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID 3</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>23.5,-22</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ,</lparam></gate>
<gate>
<ID>17</ID>
<type>AE_SMALL_INVERTER</type>
<position>96.5,-23.5</position>
<input>
<ID>IN_0</ID>135 </input>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>32,-2.5</position>
<input>
<ID>N_in1</ID>8 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>27,-9</position>
<input>
<ID>N_in0</ID>21 </input>
<input>
<ID>N_in1</ID>12 </input>
<input>
<ID>N_in3</ID>21 </input>
<gparam>LED_BOX -4.1,-1.1,4.1,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>32,-15.5</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>22,-15.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>22,-2.5</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>25</ID>
<type>GA_LED</type>
<position>27,-22</position>
<input>
<ID>N_in1</ID>15 </input>
<gparam>LED_BOX -4.1,-1.1,4.1,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>27,4</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -4.1,-1.1,4.1,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>29</ID>
<type>DE_TO</type>
<position>133,66.5</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID .</lparam></gate>
<gate>
<ID>30</ID>
<type>DE_TO</type>
<position>118,51.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>31</ID>
<type>DE_TO</type>
<position>117.5,30.5</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID '</lparam></gate>
<gate>
<ID>32</ID>
<type>DE_TO</type>
<position>117,12.5</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2</lparam></gate>
<gate>
<ID>33</ID>
<type>DE_TO</type>
<position>117,-14.5</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ,</lparam></gate>
<gate>
<ID>34</ID>
<type>DE_TO</type>
<position>114.5,0</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_AND2</type>
<position>109.5,81</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_AND2</type>
<position>109.5,77</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>DD_KEYPAD_HEX</type>
<position>48,31.5</position>
<output>
<ID>OUT_0</ID>133 </output>
<output>
<ID>OUT_1</ID>135 </output>
<output>
<ID>OUT_2</ID>134 </output>
<output>
<ID>OUT_3</ID>129 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>130</ID>
<type>AE_OR4</type>
<position>116,84</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>136 </input>
<input>
<ID>IN_2</ID>126 </input>
<input>
<ID>IN_3</ID>125 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>131</ID>
<type>DE_TO</type>
<position>122,84</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>134</ID>
<type>AE_SMALL_INVERTER</type>
<position>104.5,80</position>
<input>
<ID>IN_0</ID>135 </input>
<output>
<ID>OUT_0</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>135</ID>
<type>AE_SMALL_INVERTER</type>
<position>98.5,76</position>
<input>
<ID>IN_0</ID>133 </input>
<output>
<ID>OUT_0</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>137</ID>
<type>BM_NORX2</type>
<position>109.5,85</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_AND2</type>
<position>107,46.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>AE_OR4</type>
<position>111.5,30.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>143 </input>
<input>
<ID>IN_2</ID>145 </input>
<input>
<ID>IN_3</ID>146 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_AND2</type>
<position>104.5,33.5</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>135 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_AND2</type>
<position>104.5,29.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND2</type>
<position>104.5,25.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>149 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AE_SMALL_INVERTER</type>
<position>99.5,34.5</position>
<input>
<ID>IN_0</ID>134 </input>
<output>
<ID>OUT_0</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>152</ID>
<type>AE_SMALL_INVERTER</type>
<position>99.5,28.5</position>
<input>
<ID>IN_0</ID>133 </input>
<output>
<ID>OUT_0</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>153</ID>
<type>AE_SMALL_INVERTER</type>
<position>99.5,24.5</position>
<input>
<ID>IN_0</ID>135 </input>
<output>
<ID>OUT_0</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>155</ID>
<type>AE_OR2</type>
<position>112,12.5</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_AND2</type>
<position>106,10</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>155 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>BM_NORX2</type>
<position>106,14</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>AE_SMALL_INVERTER</type>
<position>101,9</position>
<input>
<ID>IN_0</ID>133 </input>
<output>
<ID>OUT_0</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>161</ID>
<type>AE_OR3</type>
<position>109.5,0</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>134 </input>
<input>
<ID>IN_2</ID>133 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>162</ID>
<type>AE_SMALL_INVERTER</type>
<position>104.5,2</position>
<input>
<ID>IN_0</ID>135 </input>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>163</ID>
<type>AE_OR4</type>
<position>110,-14.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<input>
<ID>IN_2</ID>18 </input>
<input>
<ID>IN_3</ID>19 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_AND2</type>
<position>101.5,-13.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>135 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_AND2</type>
<position>101,-18</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>163 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>AE_SMALL_INVERTER</type>
<position>88.5,-12.5</position>
<input>
<ID>IN_0</ID>134 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>169</ID>
<type>AE_SMALL_INVERTER</type>
<position>94,-19</position>
<input>
<ID>IN_0</ID>133 </input>
<output>
<ID>OUT_0</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>170</ID>
<type>AE_OR4</type>
<position>127,66.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>129 </input>
<input>
<ID>IN_2</ID>172 </input>
<input>
<ID>IN_3</ID>173 </input>
<output>
<ID>OUT</ID>164 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>185</ID>
<type>BM_NORX2</type>
<position>121,65.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>186</ID>
<type>AA_AND2</type>
<position>121,61.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,51.5,116,51.5</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,53.5,110,53.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-4,22,-3.5</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<connection>
<GID>8</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,46.5,110,49.5</points>
<connection>
<GID>143</GID>
<name>OUT</name></connection>
<connection>
<GID>3</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-7,32,-1.5</points>
<connection>
<GID>20</GID>
<name>N_in1</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>13</ID>
<points>25.5,4,28,4</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<connection>
<GID>9</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,50.5,110,51.5</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<connection>
<GID>7</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>25.5,-9,26,-9</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<connection>
<GID>21</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-17,22,-16.5</points>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-17,32,-16.5</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>25.5,-22,26,-22</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>25</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-11.5,105.5,-7</points>
<intersection>-11.5 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-7,105.5,-7</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-11.5,107,-11.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-13.5,107,-13.5</points>
<connection>
<GID>163</GID>
<name>IN_1</name></connection>
<connection>
<GID>166</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-18,104.5,-15.5</points>
<intersection>-18 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-15.5,107,-15.5</points>
<connection>
<GID>163</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-18,104.5,-18</points>
<connection>
<GID>167</GID>
<name>OUT</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-23.5,105.5,-17.5</points>
<intersection>-23.5 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-17.5,107,-17.5</points>
<connection>
<GID>163</GID>
<name>IN_3</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-23.5,105.5,-23.5</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-23.5,98.5,-23.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-10,27,-9</points>
<connection>
<GID>21</GID>
<name>N_in3</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-9,28,-9</points>
<connection>
<GID>21</GID>
<name>N_in0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>120,84,120,84</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<connection>
<GID>131</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,77,113,81</points>
<connection>
<GID>130</GID>
<name>IN_3</name></connection>
<intersection>77 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>112.5,77,113,77</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,81,112.5,83</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,83,113,83</points>
<connection>
<GID>130</GID>
<name>IN_2</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,36.5,55.5,88</points>
<intersection>36.5 2</intersection>
<intersection>68 6</intersection>
<intersection>88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,88,113,88</points>
<intersection>55.5 0</intersection>
<intersection>113 23</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,36.5,108.5,36.5</points>
<intersection>53 29</intersection>
<intersection>55.5 0</intersection>
<intersection>108.5 21</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>55.5,68,124,68</points>
<intersection>55.5 0</intersection>
<intersection>124 24</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>108.5,33.5,108.5,36.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>36.5 2</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>113,87,113,88</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>88 1</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>124,67.5,124,68</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>68 6</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>53,34.5,53,36.5</points>
<connection>
<GID>129</GID>
<name>OUT_3</name></connection>
<intersection>36.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,80,106.5,80</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,76,106.5,76</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,28.5,97.5,28.5</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>67.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>67.5,-25.5,67.5,84</points>
<intersection>-25.5 47</intersection>
<intersection>-19 42</intersection>
<intersection>-8 40</intersection>
<intersection>-2 22</intersection>
<intersection>9 30</intersection>
<intersection>13 18</intersection>
<intersection>28.5 1</intersection>
<intersection>45.5 37</intersection>
<intersection>60.5 28</intersection>
<intersection>64.5 38</intersection>
<intersection>76 8</intersection>
<intersection>84 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>67.5,84,106.5,84</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>67.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>67.5,76,96.5,76</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>67.5 5</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>67.5,13,103,13</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>67.5 5</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>67.5,-2,106.5,-2</points>
<connection>
<GID>161</GID>
<name>IN_2</name></connection>
<intersection>67.5 5</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>67.5,60.5,118,60.5</points>
<connection>
<GID>186</GID>
<name>IN_1</name></connection>
<intersection>67.5 5</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>67.5,9,99,9</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>67.5 5</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>67.5,45.5,104,45.5</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>67.5 5</intersection>
<intersection>71.5 44</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>67.5,64.5,118,64.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>67.5 5</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>67.5,-8,98,-8</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>67.5 5</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>67.5,-19,92,-19</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>67.5 5</intersection></hsegment>
<vsegment>
<ID>44</ID>
<points>71.5,45.5,71.5,49.5</points>
<intersection>45.5 37</intersection>
<intersection>49.5 45</intersection></vsegment>
<hsegment>
<ID>45</ID>
<points>71.5,49.5,104,49.5</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>71.5 44</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>67.5,-25.5,98.5,-25.5</points>
<connection>
<GID>13</GID>
<name>IN_2</name></connection>
<intersection>67.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-21.5,58.5,82</points>
<intersection>-21.5 41</intersection>
<intersection>-12.5 37</intersection>
<intersection>-6 35</intersection>
<intersection>0 17</intersection>
<intersection>15 30</intersection>
<intersection>26.5 15</intersection>
<intersection>34.5 5</intersection>
<intersection>53.5 39</intersection>
<intersection>62.5 25</intersection>
<intersection>66.5 11</intersection>
<intersection>78 1</intersection>
<intersection>82 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,78,106.5,78</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>58.5,82,106.5,82</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>53,34.5,97.5,34.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>53 42</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>58.5,66.5,118,66.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>58.5,26.5,101.5,26.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>58.5,0,106.5,0</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>58.5,62.5,118,62.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>58.5,15,103,15</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>58.5,-6,98,-6</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>58.5,-12.5,86.5,-12.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>58.5,53.5,106,53.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>58.5,-21.5,98.5,-21.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<vsegment>
<ID>42</ID>
<points>53,32.5,53,34.5</points>
<connection>
<GID>129</GID>
<name>OUT_2</name></connection>
<intersection>34.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-23.5,63.5,86</points>
<intersection>-23.5 33</intersection>
<intersection>-17 28</intersection>
<intersection>-14.5 18</intersection>
<intersection>2 16</intersection>
<intersection>11 25</intersection>
<intersection>24.5 12</intersection>
<intersection>30.5 1</intersection>
<intersection>32.5 8</intersection>
<intersection>47.5 26</intersection>
<intersection>51.5 31</intersection>
<intersection>69.5 22</intersection>
<intersection>80 2</intersection>
<intersection>86 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,30.5,101.5,30.5</points>
<connection>
<GID>129</GID>
<name>OUT_1</name></connection>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,80,102.5,80</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>63.5,86,106.5,86</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>63.5,32.5,101.5,32.5</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>63.5,24.5,97.5,24.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>63.5,2,102.5,2</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>63.5,-14.5,98.5,-14.5</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>63.5,69.5,124,69.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>63.5,11,103,11</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>63.5,47.5,104,47.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>63.5,-17,98,-17</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>63.5,51.5,104,51.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>63.5,-23.5,94.5,-23.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>112.5,85,113,85</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<connection>
<GID>137</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,31.5,107.5,33.5</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>31.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>107.5,31.5,108.5,31.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107.5,29.5,108.5,29.5</points>
<connection>
<GID>146</GID>
<name>IN_2</name></connection>
<connection>
<GID>148</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,25.5,108,27.5</points>
<intersection>25.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,25.5,108,25.5</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108,27.5,108.5,27.5</points>
<connection>
<GID>146</GID>
<name>IN_3</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,34.5,101.5,34.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,28.5,101.5,28.5</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,24.5,101.5,24.5</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,30.5,115.5,30.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<connection>
<GID>146</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,12.5,115,12.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<connection>
<GID>155</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,10,109,11.5</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<connection>
<GID>155</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,13.5,109,14</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<connection>
<GID>155</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,9,103,9</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,0,112.5,0</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,2,106.5,2</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114,-14.5,115,-14.5</points>
<connection>
<GID>163</GID>
<name>OUT</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-12.5,98.5,-12.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-19,98,-19</points>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection>
<connection>
<GID>167</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,66.5,131,66.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<connection>
<GID>170</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,65.5,124,65.5</points>
<connection>
<GID>170</GID>
<name>IN_2</name></connection>
<connection>
<GID>185</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,61.5,124,63.5</points>
<connection>
<GID>186</GID>
<name>OUT</name></connection>
<connection>
<GID>170</GID>
<name>IN_3</name></connection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>64.4529,-42.3596,148.472,-129.991</PageViewport>
<gate>
<ID>45</ID>
<type>GA_LED</type>
<position>99.5,-82.5</position>
<gparam>LED_BOX -30,-20,30,20</gparam>
<gparam>angle 0.0</gparam></gate></page 2>
<page 3>
<PageViewport>-12.9057,46.3721,341.152,-322.905</PageViewport></page 3>
<page 4>
<PageViewport>-12.9057,46.3721,341.152,-322.905</PageViewport></page 4>
<page 5>
<PageViewport>-12.9057,46.3721,341.152,-322.905</PageViewport></page 5>
<page 6>
<PageViewport>-12.9057,46.3721,341.152,-322.905</PageViewport></page 6>
<page 7>
<PageViewport>-12.9057,46.3721,341.152,-322.905</PageViewport></page 7>
<page 8>
<PageViewport>-12.9057,46.3721,341.152,-322.905</PageViewport></page 8>
<page 9>
<PageViewport>-12.9057,46.3721,341.152,-322.905</PageViewport></page 9></circuit>