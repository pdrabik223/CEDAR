<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-93.3168,126.735,132.984,8.74772</PageViewport>
<gate>
<ID>593</ID>
<type>GA_LED</type>
<position>2,71</position>
<input>
<ID>N_in0</ID>366 </input>
<gparam>LED_BOX -30,-20,30,20</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>594</ID>
<type>AA_TOGGLE</type>
<position>-32.5,71</position>
<output>
<ID>OUT_0</ID>366 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>CC_PULSE</type>
<position>-3.5,17</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>27</ID>
<type>CC_PULSE</type>
<position>0.5,39.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>28</ID>
<type>CC_PULSE</type>
<position>-3.5,39.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>29</ID>
<type>CC_PULSE</type>
<position>-7.5,39.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>30</ID>
<type>CC_PULSE</type>
<position>0.5,32</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>31</ID>
<type>CC_PULSE</type>
<position>-3.5,32</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>32</ID>
<type>CC_PULSE</type>
<position>-7.5,32</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>33</ID>
<type>CC_PULSE</type>
<position>0.5,24.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>34</ID>
<type>CC_PULSE</type>
<position>-3.5,24.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>35</ID>
<type>CC_PULSE</type>
<position>-7.5,24.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>-7.5,43.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>616</ID>
<type>GA_LED</type>
<position>21.5,79</position>
<input>
<ID>N_in2</ID>370 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>-3.5,43.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>617</ID>
<type>GA_LED</type>
<position>15,72.5</position>
<input>
<ID>N_in0</ID>371 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>0.5,43.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>618</ID>
<type>GA_LED</type>
<position>8.5,79</position>
<input>
<ID>N_in2</ID>367 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>-7.5,36</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>619</ID>
<type>GA_LED</type>
<position>15,85.5</position>
<input>
<ID>N_in2</ID>368 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>-3.5,36</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>620</ID>
<type>GA_LED</type>
<position>21.5,66</position>
<input>
<ID>N_in3</ID>373 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>41</ID>
<type>DE_TO</type>
<position>0.5,36</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>621</ID>
<type>GA_LED</type>
<position>8.5,66</position>
<input>
<ID>N_in0</ID>372 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>-7.5,28.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>622</ID>
<type>GA_LED</type>
<position>15,59.5</position>
<input>
<ID>N_in2</ID>374 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>-3.5,28.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>0.5,28.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>-3.5,21</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>644</ID>
<type>GA_LED</type>
<position>4,79</position>
<input>
<ID>N_in2</ID>377 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>645</ID>
<type>GA_LED</type>
<position>-2.5,72.5</position>
<input>
<ID>N_in0</ID>378 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>646</ID>
<type>GA_LED</type>
<position>-9,79</position>
<input>
<ID>N_in2</ID>375 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>647</ID>
<type>GA_LED</type>
<position>-2.5,85.5</position>
<input>
<ID>N_in2</ID>376 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>648</ID>
<type>GA_LED</type>
<position>4,66</position>
<input>
<ID>N_in3</ID>380 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>649</ID>
<type>GA_LED</type>
<position>-9,66</position>
<input>
<ID>N_in0</ID>379 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>650</ID>
<type>GA_LED</type>
<position>-2.5,59.5</position>
<input>
<ID>N_in2</ID>381 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>651</ID>
<type>DA_FROM</type>
<position>-8,97</position>
<input>
<ID>IN_0</ID>381 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b7</lparam></gate>
<gate>
<ID>652</ID>
<type>DA_FROM</type>
<position>-6,97</position>
<input>
<ID>IN_0</ID>380 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b6</lparam></gate>
<gate>
<ID>653</ID>
<type>DA_FROM</type>
<position>-4,97</position>
<input>
<ID>IN_0</ID>379 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b5</lparam></gate>
<gate>
<ID>654</ID>
<type>DA_FROM</type>
<position>-2,97</position>
<input>
<ID>IN_0</ID>378 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b4</lparam></gate>
<gate>
<ID>655</ID>
<type>DA_FROM</type>
<position>0,97</position>
<input>
<ID>IN_0</ID>377 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b3</lparam></gate>
<gate>
<ID>656</ID>
<type>DA_FROM</type>
<position>2,97</position>
<input>
<ID>IN_0</ID>376 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b2</lparam></gate>
<gate>
<ID>77</ID>
<type>CC_PULSE</type>
<position>10,17</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>657</ID>
<type>DA_FROM</type>
<position>4,97</position>
<input>
<ID>IN_0</ID>375 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b1</lparam></gate>
<gate>
<ID>78</ID>
<type>DE_TO</type>
<position>10,21</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>658</ID>
<type>GA_LED</type>
<position>-13,79</position>
<input>
<ID>N_in2</ID>384 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>659</ID>
<type>GA_LED</type>
<position>-19.5,72.5</position>
<input>
<ID>N_in0</ID>385 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>660</ID>
<type>GA_LED</type>
<position>-26,79</position>
<input>
<ID>N_in2</ID>382 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>661</ID>
<type>GA_LED</type>
<position>-19.5,85.5</position>
<input>
<ID>N_in2</ID>383 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>662</ID>
<type>GA_LED</type>
<position>-13,66</position>
<input>
<ID>N_in3</ID>387 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>663</ID>
<type>GA_LED</type>
<position>-26,66</position>
<input>
<ID>N_in0</ID>386 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>664</ID>
<type>GA_LED</type>
<position>-19.5,59.5</position>
<input>
<ID>N_in2</ID>388 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>665</ID>
<type>DA_FROM</type>
<position>-25,97</position>
<input>
<ID>IN_0</ID>388 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c7</lparam></gate>
<gate>
<ID>666</ID>
<type>DA_FROM</type>
<position>-23,97</position>
<input>
<ID>IN_0</ID>387 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c6</lparam></gate>
<gate>
<ID>667</ID>
<type>DA_FROM</type>
<position>-21,97</position>
<input>
<ID>IN_0</ID>386 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c5</lparam></gate>
<gate>
<ID>668</ID>
<type>DA_FROM</type>
<position>-19,97</position>
<input>
<ID>IN_0</ID>385 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c4</lparam></gate>
<gate>
<ID>669</ID>
<type>DA_FROM</type>
<position>-17,97</position>
<input>
<ID>IN_0</ID>384 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c3</lparam></gate>
<gate>
<ID>670</ID>
<type>DA_FROM</type>
<position>-15,97</position>
<input>
<ID>IN_0</ID>383 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c2</lparam></gate>
<gate>
<ID>671</ID>
<type>DA_FROM</type>
<position>-13,97</position>
<input>
<ID>IN_0</ID>382 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c1</lparam></gate>
<gate>
<ID>561</ID>
<type>DA_FROM</type>
<position>9.5,97</position>
<input>
<ID>IN_0</ID>374 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a7</lparam></gate>
<gate>
<ID>562</ID>
<type>DA_FROM</type>
<position>11.5,97</position>
<input>
<ID>IN_0</ID>373 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a6</lparam></gate>
<gate>
<ID>563</ID>
<type>DA_FROM</type>
<position>13.5,97</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a5</lparam></gate>
<gate>
<ID>564</ID>
<type>DA_FROM</type>
<position>15.5,97</position>
<input>
<ID>IN_0</ID>371 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a4</lparam></gate>
<gate>
<ID>571</ID>
<type>DA_FROM</type>
<position>17.5,97</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a3</lparam></gate>
<gate>
<ID>572</ID>
<type>DA_FROM</type>
<position>19.5,97</position>
<input>
<ID>IN_0</ID>368 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a2</lparam></gate>
<gate>
<ID>573</ID>
<type>DA_FROM</type>
<position>21.5,97</position>
<input>
<ID>IN_0</ID>367 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a1</lparam></gate>
<wire>
<ID>386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,65,-25,73.5</points>
<intersection>65 4</intersection>
<intersection>73.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-14,73.5,-14,95</points>
<intersection>73.5 2</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-25,73.5,-14,73.5</points>
<intersection>-25 0</intersection>
<intersection>-14 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-21,95,-14,95</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-26,65,-25,65</points>
<connection>
<GID>663</GID>
<name>N_in0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,66,-14,95</points>
<connection>
<GID>662</GID>
<name>N_in3</name></connection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-23,95,-14,95</points>
<intersection>-23 5</intersection>
<intersection>-14 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-23,95,-23,95</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<intersection>95 2</intersection></vsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,60.5,-14,95</points>
<intersection>60.5 4</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-25,95,-14,95</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-19.5,60.5,-14,60.5</points>
<connection>
<GID>664</GID>
<name>N_in2</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,41.5,-7.5,41.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,41.5,-3.5,41.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,41.5,0.5,41.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection></vsegment>
<vsegment>
<ID>2</ID>
<points>0.5,41.5,0.5,41.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,34,-7.5,34</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,34,-3.5,34</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>0.5,34,0.5,34</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<connection>
<GID>41</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,26.5,-7.5,26.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,26.5,-3.5,26.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,26.5,0.5,26.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection></vsegment>
<vsegment>
<ID>2</ID>
<points>0.5,26.5,0.5,26.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,19,-3.5,19</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,19,10,19</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-30.5,71,1,71</points>
<connection>
<GID>594</GID>
<name>OUT_0</name></connection>
<connection>
<GID>593</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,73.5,20.5,95</points>
<intersection>73.5 1</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,73.5,20.5,73.5</points>
<intersection>9.5 2</intersection>
<intersection>20.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>9.5,73.5,9.5,79</points>
<connection>
<GID>618</GID>
<name>N_in2</name></connection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>20.5,95,21.5,95</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,86.5,20.5,95</points>
<intersection>86.5 3</intersection>
<intersection>95 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>15,86.5,20.5,86.5</points>
<connection>
<GID>619</GID>
<name>N_in2</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>19.5,95,20.5,95</points>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,79,20.5,95</points>
<intersection>79 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,79,22.5,79</points>
<connection>
<GID>616</GID>
<name>N_in2</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,95,20.5,95</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,72.5,20.5,95</points>
<intersection>72.5 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,72.5,20.5,72.5</points>
<connection>
<GID>617</GID>
<name>N_in0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,95,20.5,95</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,65,9.5,71.5</points>
<intersection>65 4</intersection>
<intersection>71.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>20.5,71.5,20.5,95</points>
<intersection>71.5 2</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9.5,71.5,20.5,71.5</points>
<intersection>9.5 0</intersection>
<intersection>20.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>13.5,95,20.5,95</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<intersection>20.5 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>8.5,65,9.5,65</points>
<connection>
<GID>621</GID>
<name>N_in0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,66,20.5,95</points>
<connection>
<GID>620</GID>
<name>N_in3</name></connection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11.5,95,20.5,95</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,60.5,20.5,95</points>
<intersection>60.5 4</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>9.5,95,20.5,95</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>15,60.5,20.5,60.5</points>
<connection>
<GID>622</GID>
<name>N_in2</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,73.5,3,95</points>
<intersection>73.5 1</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,73.5,3,73.5</points>
<intersection>-8 2</intersection>
<intersection>3 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-8,73.5,-8,79</points>
<connection>
<GID>646</GID>
<name>N_in2</name></connection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>3,95,4,95</points>
<intersection>3 0</intersection>
<intersection>4 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>4,95,4,95</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>95 3</intersection></vsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,86.5,3,95</points>
<intersection>86.5 3</intersection>
<intersection>95 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2.5,86.5,3,86.5</points>
<connection>
<GID>647</GID>
<name>N_in2</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>2,95,3,95</points>
<intersection>2 7</intersection>
<intersection>3 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>2,95,2,95</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>95 4</intersection></vsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,79,3,95</points>
<intersection>79 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,79,5,79</points>
<connection>
<GID>644</GID>
<name>N_in2</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.30078e-008,95,3,95</points>
<intersection>-7.30078e-008 4</intersection>
<intersection>3 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-7.30078e-008,95,-7.30078e-008,95</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>95 2</intersection></vsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,72.5,3,95</points>
<intersection>72.5 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,72.5,3,72.5</points>
<connection>
<GID>645</GID>
<name>N_in0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,95,3,95</points>
<intersection>-2 4</intersection>
<intersection>3 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-2,95,-2,95</points>
<connection>
<GID>654</GID>
<name>IN_0</name></connection>
<intersection>95 2</intersection></vsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,65,-8,73.5</points>
<intersection>65 4</intersection>
<intersection>73.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>3,73.5,3,95</points>
<intersection>73.5 2</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8,73.5,3,73.5</points>
<intersection>-8 0</intersection>
<intersection>3 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4,95,3,95</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>3 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-9,65,-8,65</points>
<connection>
<GID>649</GID>
<name>N_in0</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,66,3,95</points>
<connection>
<GID>648</GID>
<name>N_in3</name></connection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-6,95,3,95</points>
<intersection>-6 5</intersection>
<intersection>3 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-6,95,-6,95</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>95 2</intersection></vsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,60.5,3,95</points>
<intersection>60.5 4</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-8,95,3,95</points>
<intersection>-8 7</intersection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-2.5,60.5,3,60.5</points>
<connection>
<GID>650</GID>
<name>N_in2</name></connection>
<intersection>3 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-8,95,-8,95</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>95 3</intersection></vsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,73.5,-14,95</points>
<intersection>73.5 1</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,73.5,-14,73.5</points>
<intersection>-25 2</intersection>
<intersection>-14 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-25,73.5,-25,79</points>
<connection>
<GID>660</GID>
<name>N_in2</name></connection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-14,95,-13,95</points>
<intersection>-14 0</intersection>
<intersection>-13 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-13,95,-13,95</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>95 3</intersection></vsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,86.5,-14,95</points>
<intersection>86.5 3</intersection>
<intersection>95 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,86.5,-14,86.5</points>
<connection>
<GID>661</GID>
<name>N_in2</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-15,95,-14,95</points>
<intersection>-15 7</intersection>
<intersection>-14 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-15,95,-15,95</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>95 4</intersection></vsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,79,-14,95</points>
<intersection>79 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,79,-12,79</points>
<connection>
<GID>658</GID>
<name>N_in2</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-17,95,-14,95</points>
<intersection>-17 4</intersection>
<intersection>-14 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-17,95,-17,95</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>95 2</intersection></vsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,72.5,-14,95</points>
<intersection>72.5 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-18.5,72.5,-14,72.5</points>
<connection>
<GID>659</GID>
<name>N_in0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19,95,-14,95</points>
<intersection>-19 4</intersection>
<intersection>-14 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-19,95,-19,95</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>95 2</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-76.2543,90.493,376.347,-145.481</PageViewport>
<gate>
<ID>1</ID>
<type>BM_NORX2</type>
<position>285,29</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_OR3</type>
<position>287,65</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>3 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_SMALL_INVERTER</type>
<position>282,67</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>BM_NORX2</type>
<position>281,64</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,56</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND3</type>
<position>285,16</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>26 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,50</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,46</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_OR2</type>
<position>291,42</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>285,39</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>BM_NORX2</type>
<position>285,43</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,38</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_OR3</type>
<position>285,34</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>27 </input>
<input>
<ID>IN_2</ID>26 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,36</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>15</ID>
<type>AE_OR4</type>
<position>292,24</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>285,25</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_AND2</type>
<position>285,21</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,26</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,20</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_OR4</type>
<position>286.5,75</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>23 </input>
<input>
<ID>IN_2</ID>71 </input>
<input>
<ID>IN_3</ID>72 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>21</ID>
<type>BM_NORX2</type>
<position>280.5,74</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>280.5,70</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,16</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>285,47</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>DE_TO</type>
<position>292.5,75</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a2</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>292,65</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a3</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>298,52</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a4</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>296,42</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a5</lparam></gate>
<gate>
<ID>49</ID>
<type>DE_TO</type>
<position>298,24</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a7</lparam></gate>
<gate>
<ID>50</ID>
<type>DE_TO</type>
<position>290,34</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a6</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_AND2</type>
<position>285,85</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND2</type>
<position>285,81</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_OR4</type>
<position>291.5,88</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>29 </input>
<input>
<ID>IN_2</ID>22 </input>
<input>
<ID>IN_3</ID>21 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>54</ID>
<type>DE_TO</type>
<position>297.5,88</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a1</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,84</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>65</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>44,-23.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>41 </input>
<input>
<ID>IN_3</ID>40 </input>
<output>
<ID>OUT_0</ID>59 </output>
<output>
<ID>OUT_1</ID>55 </output>
<output>
<ID>OUT_2</ID>54 </output>
<output>
<ID>OUT_3</ID>53 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>66</ID>
<type>DE_OR8</type>
<position>31.5,-34.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>35 </input>
<input>
<ID>IN_3</ID>34 </input>
<input>
<ID>IN_4</ID>30 </input>
<input>
<ID>IN_5</ID>31 </input>
<input>
<ID>IN_6</ID>32 </input>
<input>
<ID>IN_7</ID>33 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>67</ID>
<type>FF_GND</type>
<position>27.5,-33</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_OR2</type>
<position>31.5,-12.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_OR4</type>
<position>31.5,-26.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>31 </input>
<input>
<ID>IN_3</ID>38 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>70</ID>
<type>AE_OR4</type>
<position>31.5,-18.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>32 </input>
<input>
<ID>IN_3</ID>43 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_OR4</type>
<position>45,-11.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>37 </input>
<input>
<ID>IN_3</ID>36 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_OR2</type>
<position>53,-3.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>BB_CLOCK</type>
<position>46,-46</position>
<output>
<ID>CLK</ID>61 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>52.5,-44</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_REGISTER4</type>
<position>52.5,-31.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>54 </input>
<input>
<ID>IN_3</ID>53 </input>
<input>
<ID>clear</ID>107 </input>
<input>
<ID>clock</ID>61 </input>
<input>
<ID>load</ID>58 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>79</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,80</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>80</ID>
<type>BM_NORX2</type>
<position>285,89</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_AND2</type>
<position>281,60</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AE_OR4</type>
<position>292,52</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>44 </input>
<input>
<ID>IN_2</ID>46 </input>
<input>
<ID>IN_3</ID>47 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_AND2</type>
<position>285,55</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_AND2</type>
<position>285,51</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>HA_JUNC_2</type>
<position>259,53</position>
<input>
<ID>N_in0</ID>111 </input>
<input>
<ID>N_in1</ID>26 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>HA_JUNC_2</type>
<position>259,54</position>
<input>
<ID>N_in0</ID>112 </input>
<input>
<ID>N_in1</ID>28 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>HA_JUNC_2</type>
<position>259,55</position>
<input>
<ID>N_in0</ID>113 </input>
<input>
<ID>N_in1</ID>27 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>HA_JUNC_2</type>
<position>259,56</position>
<input>
<ID>N_in0</ID>114 </input>
<input>
<ID>N_in1</ID>23 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>CC_PULSE</type>
<position>-4,-7</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>90</ID>
<type>CC_PULSE</type>
<position>0,15.5</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>91</ID>
<type>CC_PULSE</type>
<position>-4,15.5</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>92</ID>
<type>CC_PULSE</type>
<position>-8,15.5</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>93</ID>
<type>CC_PULSE</type>
<position>0,8</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>94</ID>
<type>CC_PULSE</type>
<position>-4,8</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>95</ID>
<type>CC_PULSE</type>
<position>-8,8</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>96</ID>
<type>CC_PULSE</type>
<position>0,0.5</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>97</ID>
<type>CC_PULSE</type>
<position>-4,0.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>98</ID>
<type>CC_PULSE</type>
<position>-8,0.5</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>99</ID>
<type>DE_TO</type>
<position>-8,19.5</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t7</lparam></gate>
<gate>
<ID>100</ID>
<type>DE_TO</type>
<position>-4,19.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t8</lparam></gate>
<gate>
<ID>101</ID>
<type>DE_TO</type>
<position>0,19.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t9</lparam></gate>
<gate>
<ID>102</ID>
<type>DE_TO</type>
<position>-8,12</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t4</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>-4,12</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t5</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>0,12</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t6</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>-8,4.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t1</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>-4,4.5</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t2</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_TO</type>
<position>0,4.5</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t3</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>-4,-3</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t0</lparam></gate>
<gate>
<ID>109</ID>
<type>CC_PULSE</type>
<position>-12,-10</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>-12,-6</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID tCE</lparam></gate>
<gate>
<ID>112</ID>
<type>AE_OR2</type>
<position>12,-6</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AE_OR2</type>
<position>12,-10</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_OR2</type>
<position>12,-14</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>102 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AE_OR2</type>
<position>12,-18</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>AE_OR2</type>
<position>12,-22</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_OR2</type>
<position>12,-26</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR2</type>
<position>12,-30</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>98 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_OR2</type>
<position>12,-34</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_OR2</type>
<position>12,-38</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_OR2</type>
<position>12,-42</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>7,-43</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t0</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>7,-37</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t1</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>7,-33</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t2</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>7,-29</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t3</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>7,-25</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t4</lparam></gate>
<gate>
<ID>129</ID>
<type>DA_FROM</type>
<position>7,-21</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t5</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>7,-17</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t6</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>7,-13</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t7</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>7,-9</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t8</lparam></gate>
<gate>
<ID>133</ID>
<type>DA_FROM</type>
<position>7,-5</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t9</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>7,-41</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>7,-39</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>7,-35</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>137</ID>
<type>DA_FROM</type>
<position>7,-31</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>138</ID>
<type>DA_FROM</type>
<position>7,-27</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>139</ID>
<type>DA_FROM</type>
<position>7,-23</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>140</ID>
<type>DA_FROM</type>
<position>7,-19</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>141</ID>
<type>DA_FROM</type>
<position>7,-15</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>7,-11</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>7,-7</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>144</ID>
<type>DA_FROM</type>
<position>54.5,-44</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID tCE</lparam></gate>
<gate>
<ID>145</ID>
<type>AE_OR2</type>
<position>53.5,-39</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>GA_LED</type>
<position>249.5,-9</position>
<input>
<ID>N_in0</ID>221 </input>
<input>
<ID>N_in1</ID>111 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>249.5,-12</position>
<input>
<ID>N_in0</ID>222 </input>
<input>
<ID>N_in1</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>249.5,-15</position>
<input>
<ID>N_in0</ID>223 </input>
<input>
<ID>N_in1</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>GA_LED</type>
<position>249.5,-18</position>
<input>
<ID>N_in0</ID>224 </input>
<input>
<ID>N_in1</ID>114 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>GA_LED</type>
<position>249.5,-23</position>
<input>
<ID>N_in0</ID>392 </input>
<input>
<ID>N_in1</ID>191 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>GA_LED</type>
<position>249.5,-26</position>
<input>
<ID>N_in0</ID>391 </input>
<input>
<ID>N_in1</ID>192 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>GA_LED</type>
<position>249.5,-29</position>
<input>
<ID>N_in0</ID>390 </input>
<input>
<ID>N_in1</ID>193 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>249.5,-32</position>
<input>
<ID>N_in0</ID>389 </input>
<input>
<ID>N_in1</ID>194 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>GA_LED</type>
<position>249.5,-36</position>
<input>
<ID>N_in0</ID>396 </input>
<input>
<ID>N_in1</ID>195 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>249.5,-39</position>
<input>
<ID>N_in0</ID>395 </input>
<input>
<ID>N_in1</ID>196 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>GA_LED</type>
<position>249.5,-42</position>
<input>
<ID>N_in0</ID>394 </input>
<input>
<ID>N_in1</ID>197 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>249.5,-45</position>
<input>
<ID>N_in0</ID>393 </input>
<input>
<ID>N_in1</ID>198 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>DD_KEYPAD_HEX</type>
<position>230.5,-15</position>
<output>
<ID>OUT_0</ID>221 </output>
<output>
<ID>OUT_1</ID>222 </output>
<output>
<ID>OUT_2</ID>223 </output>
<output>
<ID>OUT_3</ID>224 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 10</lparam></gate>
<gate>
<ID>161</ID>
<type>BM_NORX2</type>
<position>287,-51</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>AE_OR3</type>
<position>289,-15</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>118 </input>
<input>
<ID>IN_2</ID>117 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>163</ID>
<type>AE_SMALL_INVERTER</type>
<position>284,-13</position>
<input>
<ID>IN_0</ID>131 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>164</ID>
<type>BM_NORX2</type>
<position>283,-16</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>AE_SMALL_INVERTER</type>
<position>282,-24</position>
<input>
<ID>IN_0</ID>131 </input>
<output>
<ID>OUT_0</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_AND3</type>
<position>287,-64</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>123 </input>
<input>
<ID>IN_2</ID>130 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>167</ID>
<type>AE_SMALL_INVERTER</type>
<position>282,-30</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>168</ID>
<type>AE_SMALL_INVERTER</type>
<position>282,-34</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>169</ID>
<type>AE_OR2</type>
<position>293,-38</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND2</type>
<position>287,-41</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>BM_NORX2</type>
<position>287,-37</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AE_SMALL_INVERTER</type>
<position>282,-42</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>173</ID>
<type>AE_OR3</type>
<position>287,-46</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>131 </input>
<input>
<ID>IN_2</ID>130 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>174</ID>
<type>AE_SMALL_INVERTER</type>
<position>282,-44</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>175</ID>
<type>AE_OR4</type>
<position>294,-56</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>120 </input>
<input>
<ID>IN_2</ID>121 </input>
<input>
<ID>IN_3</ID>122 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_AND2</type>
<position>287,-55</position>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_AND2</type>
<position>287,-59</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>149 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>AE_SMALL_INVERTER</type>
<position>282,-54</position>
<input>
<ID>IN_0</ID>131 </input>
<output>
<ID>OUT_0</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>179</ID>
<type>AE_SMALL_INVERTER</type>
<position>282,-60</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>180</ID>
<type>AE_OR4</type>
<position>288.5,-5</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>127 </input>
<input>
<ID>IN_2</ID>151 </input>
<input>
<ID>IN_3</ID>152 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>181</ID>
<type>BM_NORX2</type>
<position>282.5,-6</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_AND2</type>
<position>282.5,-10</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>AE_SMALL_INVERTER</type>
<position>282,-64</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_AND2</type>
<position>287,-33</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>139 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>185</ID>
<type>DE_TO</type>
<position>294.5,-5</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b2</lparam></gate>
<gate>
<ID>186</ID>
<type>DE_TO</type>
<position>294,-15</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b3</lparam></gate>
<gate>
<ID>187</ID>
<type>DE_TO</type>
<position>300,-28</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b4</lparam></gate>
<gate>
<ID>188</ID>
<type>DE_TO</type>
<position>298,-38</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b5</lparam></gate>
<gate>
<ID>189</ID>
<type>DE_TO</type>
<position>300,-56</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b7</lparam></gate>
<gate>
<ID>190</ID>
<type>DE_TO</type>
<position>292,-46</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b6</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_AND2</type>
<position>287,5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_AND2</type>
<position>287,1</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>193</ID>
<type>AE_OR4</type>
<position>293.5,8</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>133 </input>
<input>
<ID>IN_2</ID>126 </input>
<input>
<ID>IN_3</ID>125 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>194</ID>
<type>DE_TO</type>
<position>299.5,8</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b1</lparam></gate>
<gate>
<ID>195</ID>
<type>AE_SMALL_INVERTER</type>
<position>282,4</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>196</ID>
<type>AE_SMALL_INVERTER</type>
<position>282,0</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>197</ID>
<type>BM_NORX2</type>
<position>287,9</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND2</type>
<position>283,-20</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_OR4</type>
<position>294,-28</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>134 </input>
<input>
<ID>IN_2</ID>135 </input>
<input>
<ID>IN_3</ID>136 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_AND2</type>
<position>287,-25</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_AND2</type>
<position>287,-29</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>HA_JUNC_2</type>
<position>261,-27</position>
<input>
<ID>N_in0</ID>191 </input>
<input>
<ID>N_in1</ID>130 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>HA_JUNC_2</type>
<position>261,-26</position>
<input>
<ID>N_in0</ID>192 </input>
<input>
<ID>N_in1</ID>132 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>204</ID>
<type>HA_JUNC_2</type>
<position>261,-25</position>
<input>
<ID>N_in0</ID>193 </input>
<input>
<ID>N_in1</ID>131 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>HA_JUNC_2</type>
<position>261,-24</position>
<input>
<ID>N_in0</ID>194 </input>
<input>
<ID>N_in1</ID>127 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>BM_NORX2</type>
<position>287.5,-133.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>AE_OR3</type>
<position>289.5,-97.5</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>156 </input>
<input>
<ID>IN_2</ID>155 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>208</ID>
<type>AE_SMALL_INVERTER</type>
<position>284.5,-95.5</position>
<input>
<ID>IN_0</ID>169 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>209</ID>
<type>BM_NORX2</type>
<position>283.5,-98.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>AE_SMALL_INVERTER</type>
<position>282.5,-106.5</position>
<input>
<ID>IN_0</ID>169 </input>
<output>
<ID>OUT_0</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_AND3</type>
<position>287.5,-146.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>161 </input>
<input>
<ID>IN_2</ID>168 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>212</ID>
<type>AE_SMALL_INVERTER</type>
<position>282.5,-112.5</position>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>213</ID>
<type>AE_SMALL_INVERTER</type>
<position>282.5,-116.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>214</ID>
<type>AE_OR2</type>
<position>293.5,-120.5</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>180 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_AND2</type>
<position>287.5,-123.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>182 </input>
<output>
<ID>OUT</ID>180 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>BM_NORX2</type>
<position>287.5,-119.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>AE_SMALL_INVERTER</type>
<position>282.5,-124.5</position>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>182 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>218</ID>
<type>AE_OR3</type>
<position>287.5,-128.5</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>169 </input>
<input>
<ID>IN_2</ID>168 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>219</ID>
<type>AE_SMALL_INVERTER</type>
<position>282.5,-126.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>184 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>220</ID>
<type>AE_OR4</type>
<position>294.5,-138.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>158 </input>
<input>
<ID>IN_2</ID>159 </input>
<input>
<ID>IN_3</ID>160 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>287.5,-137.5</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_AND2</type>
<position>287.5,-141.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>223</ID>
<type>AE_SMALL_INVERTER</type>
<position>282.5,-136.5</position>
<input>
<ID>IN_0</ID>169 </input>
<output>
<ID>OUT_0</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>224</ID>
<type>AE_SMALL_INVERTER</type>
<position>282.5,-142.5</position>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>225</ID>
<type>AE_OR4</type>
<position>289,-87.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>165 </input>
<input>
<ID>IN_2</ID>189 </input>
<input>
<ID>IN_3</ID>190 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>226</ID>
<type>BM_NORX2</type>
<position>283,-88.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_AND2</type>
<position>283,-92.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AE_SMALL_INVERTER</type>
<position>282.5,-146.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_AND2</type>
<position>287.5,-115.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>177 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>DE_TO</type>
<position>295.5,-87.5</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c2</lparam></gate>
<gate>
<ID>231</ID>
<type>DE_TO</type>
<position>294.5,-97.5</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c3</lparam></gate>
<gate>
<ID>232</ID>
<type>DE_TO</type>
<position>300.5,-110.5</position>
<input>
<ID>IN_0</ID>178 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c4</lparam></gate>
<gate>
<ID>233</ID>
<type>DE_TO</type>
<position>298.5,-120.5</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c5</lparam></gate>
<gate>
<ID>234</ID>
<type>DE_TO</type>
<position>300.5,-138.5</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c7</lparam></gate>
<gate>
<ID>235</ID>
<type>DE_TO</type>
<position>292.5,-128.5</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c6</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>287.5,-77.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>166 </input>
<output>
<ID>OUT</ID>164 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>AA_AND2</type>
<position>287.5,-81.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>167 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>238</ID>
<type>AE_OR4</type>
<position>294,-74.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>171 </input>
<input>
<ID>IN_2</ID>164 </input>
<input>
<ID>IN_3</ID>163 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>239</ID>
<type>DE_TO</type>
<position>300,-74.5</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c1</lparam></gate>
<gate>
<ID>240</ID>
<type>AE_SMALL_INVERTER</type>
<position>282.5,-78.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_SMALL_INVERTER</type>
<position>282.5,-82.5</position>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>167 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>242</ID>
<type>BM_NORX2</type>
<position>287.5,-73.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_AND2</type>
<position>283.5,-102.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>AE_OR4</type>
<position>294.5,-110.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>172 </input>
<input>
<ID>IN_2</ID>173 </input>
<input>
<ID>IN_3</ID>174 </input>
<output>
<ID>OUT</ID>178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>245</ID>
<type>AA_AND2</type>
<position>287.5,-107.5</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_AND2</type>
<position>287.5,-111.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>176 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>247</ID>
<type>HA_JUNC_2</type>
<position>261.5,-109.5</position>
<input>
<ID>N_in0</ID>195 </input>
<input>
<ID>N_in1</ID>168 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>HA_JUNC_2</type>
<position>261.5,-108.5</position>
<input>
<ID>N_in0</ID>196 </input>
<input>
<ID>N_in1</ID>170 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>249</ID>
<type>HA_JUNC_2</type>
<position>261.5,-107.5</position>
<input>
<ID>N_in0</ID>197 </input>
<input>
<ID>N_in1</ID>169 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>HA_JUNC_2</type>
<position>261.5,-106.5</position>
<input>
<ID>N_in0</ID>198 </input>
<input>
<ID>N_in1</ID>165 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>672</ID>
<type>DD_KEYPAD_HEX</type>
<position>230.5,-27</position>
<output>
<ID>OUT_0</ID>392 </output>
<output>
<ID>OUT_1</ID>391 </output>
<output>
<ID>OUT_2</ID>390 </output>
<output>
<ID>OUT_3</ID>389 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 8</lparam></gate>
<gate>
<ID>673</ID>
<type>DD_KEYPAD_HEX</type>
<position>230,-39</position>
<output>
<ID>OUT_0</ID>396 </output>
<output>
<ID>OUT_1</ID>395 </output>
<output>
<ID>OUT_2</ID>394 </output>
<output>
<ID>OUT_3</ID>393 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-32,242,-24</points>
<intersection>-32 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242,-32,248.5,-32</points>
<connection>
<GID>154</GID>
<name>N_in0</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235.5,-24,242,-24</points>
<connection>
<GID>672</GID>
<name>OUT_3</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-29,242,-26</points>
<intersection>-29 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242,-29,248.5,-29</points>
<connection>
<GID>153</GID>
<name>N_in0</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235.5,-26,242,-26</points>
<connection>
<GID>672</GID>
<name>OUT_2</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,65,290,65</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-28,242,-26</points>
<intersection>-28 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242,-26,248.5,-26</points>
<connection>
<GID>152</GID>
<name>N_in0</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235.5,-28,242,-28</points>
<connection>
<GID>672</GID>
<name>OUT_1</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,67,284,67</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-30,242,-23</points>
<intersection>-30 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235.5,-30,242,-30</points>
<connection>
<GID>672</GID>
<name>OUT_0</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242,-23,248.5,-23</points>
<connection>
<GID>151</GID>
<name>N_in0</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,60,284,63</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-45,241.5,-36</points>
<intersection>-45 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241.5,-45,248.5,-45</points>
<connection>
<GID>158</GID>
<name>N_in0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235,-36,241.5,-36</points>
<connection>
<GID>673</GID>
<name>OUT_3</name></connection>
<intersection>241.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-42,241.5,-38</points>
<intersection>-42 2</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,-38,241.5,-38</points>
<connection>
<GID>673</GID>
<name>OUT_2</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>241.5,-42,248.5,-42</points>
<connection>
<GID>157</GID>
<name>N_in0</name></connection>
<intersection>241.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-40,241.5,-39</points>
<intersection>-40 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241.5,-39,248.5,-39</points>
<connection>
<GID>156</GID>
<name>N_in0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235,-40,241.5,-40</points>
<connection>
<GID>673</GID>
<name>OUT_1</name></connection>
<intersection>241.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-42,241.5,-36</points>
<intersection>-42 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,-42,241.5,-42</points>
<connection>
<GID>673</GID>
<name>OUT_0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>241.5,-36,248.5,-36</points>
<connection>
<GID>155</GID>
<name>N_in0</name></connection>
<intersection>241.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,64,284,65</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,27,289,29</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288,29,289,29</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288,25,289,25</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<connection>
<GID>16</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,21,288,23</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288,23,289,23</points>
<connection>
<GID>15</GID>
<name>IN_2</name></connection>
<intersection>288 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,16,289,21</points>
<connection>
<GID>15</GID>
<name>IN_3</name></connection>
<intersection>16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>288,16,289,16</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,16,282,16</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,88,295.5,88</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<connection>
<GID>54</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,81,288.5,85</points>
<connection>
<GID>53</GID>
<name>IN_3</name></connection>
<intersection>81 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>288,81,288.5,81</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,85,288,87</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288,87,288.5,87</points>
<connection>
<GID>53</GID>
<name>IN_2</name></connection>
<intersection>288 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266,56,266,91</points>
<intersection>56 2</intersection>
<intersection>76 6</intersection>
<intersection>91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,91,288.5,91</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>266 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>260,56,289,56</points>
<connection>
<GID>88</GID>
<name>N_in1</name></connection>
<intersection>266 0</intersection>
<intersection>289 21</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>266,76,283.5,76</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>266 0</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>289,55,289,56</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>56 2</intersection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,84,282,84</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>282,80,282,80</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>265.5,50,278,50</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>265.5 50</intersection>
<intersection>278 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>278,14,278,88</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>14 47</intersection>
<intersection>28 40</intersection>
<intersection>32 22</intersection>
<intersection>42 18</intersection>
<intersection>50 1</intersection>
<intersection>69 28</intersection>
<intersection>73 38</intersection>
<intersection>88 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>278,88,282,88</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>278 5</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>278,42,282,42</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>278 5</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>278,32,282,32</points>
<connection>
<GID>13</GID>
<name>IN_2</name></connection>
<intersection>278 5</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>277.5,69,278,69</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>278 5</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>277.5,73,278,73</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>278 5</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>278,28,282,28</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>278 5</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>278,14,282,14</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>278 5</intersection></hsegment>
<vsegment>
<ID>50</ID>
<points>265.5,50,265.5,53</points>
<intersection>50 1</intersection>
<intersection>53 51</intersection></vsegment>
<hsegment>
<ID>51</ID>
<points>260,53,265.5,53</points>
<connection>
<GID>85</GID>
<name>N_in1</name></connection>
<intersection>265.5 50</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,18,269,86</points>
<intersection>18 41</intersection>
<intersection>26 37</intersection>
<intersection>30 35</intersection>
<intersection>34 17</intersection>
<intersection>44 30</intersection>
<intersection>48 15</intersection>
<intersection>55 45</intersection>
<intersection>56 5</intersection>
<intersection>67 39</intersection>
<intersection>71 25</intersection>
<intersection>75 11</intersection>
<intersection>82 1</intersection>
<intersection>86 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269,82,282,82</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>269,86,282,86</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>269,56,278,56</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>269,75,277.5,75</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>269,48,282,48</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>269,34,282,34</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>269,71,277.5,71</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>269,44,282,44</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>269,30,282,30</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>269,26,278,26</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>269,67,280,67</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>269,18,282,18</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>260,55,269,55</points>
<connection>
<GID>87</GID>
<name>N_in1</name></connection>
<intersection>269 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,16,274,90</points>
<intersection>16 33</intersection>
<intersection>22 28</intersection>
<intersection>24 18</intersection>
<intersection>36 16</intersection>
<intersection>40 25</intersection>
<intersection>46 12</intersection>
<intersection>54 8</intersection>
<intersection>61 26</intersection>
<intersection>65 31</intersection>
<intersection>78 1</intersection>
<intersection>84 2</intersection>
<intersection>90 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264.5,78,283.5,78</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>264.5 36</intersection>
<intersection>274 0</intersection>
<intersection>282 38</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274,84,278,84</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>274,90,282,90</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>260,54,282,54</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<connection>
<GID>86</GID>
<name>N_in1</name></connection>
<intersection>264.5 36</intersection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>274,46,278,46</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>274,36,278,36</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>274,24,282,24</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>274,40,282,40</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>274,61,278,61</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>274,22,282,22</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>274,65,278,65</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>274,16,278,16</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>274 0</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>264.5,54,264.5,78</points>
<intersection>54 8</intersection>
<intersection>78 1</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>282,52,282,78</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>78 1</intersection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288,89,288.5,89</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<connection>
<GID>80</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>15,-38,28.5,-38</points>
<connection>
<GID>66</GID>
<name>IN_4</name></connection>
<connection>
<GID>120</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-37,24,-27.5</points>
<intersection>-37 2</intersection>
<intersection>-30 4</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24,-37,28.5,-37</points>
<connection>
<GID>66</GID>
<name>IN_5</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24,-27.5,28.5,-27.5</points>
<connection>
<GID>69</GID>
<name>IN_2</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>15,-30,24,-30</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-36,24.5,-19.5</points>
<intersection>-36 2</intersection>
<intersection>-22.5 1</intersection>
<intersection>-19.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-22.5,24.5,-22.5</points>
<intersection>15 4</intersection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-36,28.5,-36</points>
<connection>
<GID>66</GID>
<name>IN_6</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24.5,-19.5,28.5,-19.5</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>24.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-22.5,15,-22</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>-22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-35,25,-15.5</points>
<intersection>-35 2</intersection>
<intersection>-23.5 3</intersection>
<intersection>-18.5 1</intersection>
<intersection>-15.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-18.5,25,-18.5</points>
<intersection>15 5</intersection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-35,28.5,-35</points>
<connection>
<GID>66</GID>
<name>IN_7</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25,-23.5,28.5,-23.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>25,-15.5,28.5,-15.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>15,-18.5,15,-14</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-34,25.5,-6</points>
<intersection>-34 2</intersection>
<intersection>-11.5 3</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-6,25.5,-6</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-34,28.5,-34</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25.5,-11.5,28.5,-11.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-33,28.5,-31</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-34.5,37,-14.5</points>
<intersection>-34.5 8</intersection>
<intersection>-24.5 4</intersection>
<intersection>-14.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37,-24.5,41,-24.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>37,-14.5,42,-14.5</points>
<connection>
<GID>72</GID>
<name>IN_3</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>35.5,-34.5,37,-34.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-26.5,36.5,-12.5</points>
<intersection>-26.5 2</intersection>
<intersection>-23.5 1</intersection>
<intersection>-12.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-23.5,41,-23.5</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-26.5,36.5,-26.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36.5,-12.5,42,-12.5</points>
<connection>
<GID>72</GID>
<name>IN_2</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-29.5,24,-28.5</points>
<intersection>-29.5 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-28.5,24,-28.5</points>
<intersection>20.5 3</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-29.5,28.5,-29.5</points>
<connection>
<GID>69</GID>
<name>IN_3</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20.5,-34,20.5,-28.5</points>
<intersection>-34 4</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>15,-34,20.5,-34</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>20.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-25.5,24,-17.5</points>
<intersection>-25.5 2</intersection>
<intersection>-20.5 1</intersection>
<intersection>-17.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-20.5,24,-20.5</points>
<intersection>15 4</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-25.5,28.5,-25.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24,-17.5,28.5,-17.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-20.5,15,-18</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-21.5,38,-12.5</points>
<intersection>-21.5 3</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-12.5,38,-12.5</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38,-21.5,41,-21.5</points>
<connection>
<GID>65</GID>
<name>IN_3</name></connection>
<intersection>38 0</intersection>
<intersection>40 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>40,-21.5,40,-8.5</points>
<intersection>-21.5 3</intersection>
<intersection>-8.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>40,-8.5,42,-8.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>40 6</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-22.5,36.5,-18.5</points>
<intersection>-22.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-22.5,41,-22.5</points>
<connection>
<GID>65</GID>
<name>IN_2</name></connection>
<intersection>36.5 0</intersection>
<intersection>39 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-18.5,36.5,-18.5</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>39,-22.5,39,-10.5</points>
<intersection>-22.5 1</intersection>
<intersection>-10.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>39,-10.5,42,-10.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>39 5</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-16.5,24.5,-13.5</points>
<intersection>-16.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-16.5,24.5,-16.5</points>
<intersection>15 3</intersection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-13.5,28.5,-13.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,-16.5,15,-10</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>-16.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-24.5,24,-21.5</points>
<intersection>-24.5 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-24.5,24,-24.5</points>
<intersection>15 3</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-21.5,28.5,-21.5</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,-26,15,-24.5</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,53,288,55</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>288,53,289,53</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>288 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-42,22,-4.5</points>
<intersection>-42 4</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22,-4.5,50,-4.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>15,-42,22,-42</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288,51,289,51</points>
<connection>
<GID>82</GID>
<name>IN_2</name></connection>
<connection>
<GID>84</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,47,288.5,49</points>
<intersection>47 1</intersection>
<intersection>49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288,47,288.5,47</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>288.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>288.5,49,289,49</points>
<connection>
<GID>82</GID>
<name>IN_3</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,56,282,56</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<connection>
<GID>83</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,50,282,50</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,46,282,46</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296,52,296,52</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>82</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,42,294,42</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-29.5,42.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_3</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-29.5,48.5,-29.5</points>
<connection>
<GID>76</GID>
<name>IN_3</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-30.5,43.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_2</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-30.5,48.5,-30.5</points>
<connection>
<GID>76</GID>
<name>IN_2</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-31.5,44.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_1</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-31.5,48.5,-31.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,39,288,41</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<connection>
<GID>9</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-11.5,49,-2.5</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-2.5,50,-2.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-26.5,51.5,-15.5</points>
<connection>
<GID>76</GID>
<name>load</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-15.5,56,-15.5</points>
<intersection>51.5 0</intersection>
<intersection>56 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>56,-15.5,56,-3.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>-15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-32.5,45.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-32.5,48.5,-32.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-42,46,-35.5</points>
<connection>
<GID>74</GID>
<name>CLK</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-35.5,51.5,-35.5</points>
<connection>
<GID>76</GID>
<name>clock</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,43,288,43</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>11</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,38,282,38</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,34,288,34</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<connection>
<GID>50</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,36,282,36</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296,24,296,24</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<connection>
<GID>49</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,26,282,26</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,20,282,20</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,75,290.5,75</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>283.5,74,283.5,74</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<connection>
<GID>21</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>283.5,70,283.5,72</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-8,17.5,-8,17.5</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,17.5,-4,17.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>17.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-4,17.5,-4,17.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.43359e-008,17.5,2.43359e-008,17.5</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection></vsegment>
<vsegment>
<ID>2</ID>
<points>-2.43359e-008,17.5,-2.43359e-008,17.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,10,-8,10</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>10 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-8,10,-8,10</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,10,-4,10</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>10 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-4,10,-4,10</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-2.43359e-008,10,2.43359e-008,10</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>-2.43359e-008 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>-2.43359e-008,10,-2.43359e-008,10</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>10 0</intersection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,2.5,-8,2.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>2.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-8,2.5,-8,2.5</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,2.5,-4,2.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>2.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-4,2.5,-4,2.5</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.43359e-008,2.5,2.43359e-008,2.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection></vsegment>
<vsegment>
<ID>2</ID>
<points>-2.43359e-008,2.5,-2.43359e-008,2.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-5,-4,-5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-4,-5,-4,-5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-8,-12,-8</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>-8 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-12,-8,-12,-8</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-43,9,-43</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-43,9,-43</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-37,9,-37</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-37,9,-37</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-33,9,-33</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-33,9,-33</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-29,9,-29</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-29,9,-29</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-25,9,-25</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-25,9,-25</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-21,9,-21</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-21,9,-21</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-17,9,-17</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-17,9,-17</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-13,9,-13</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-13,9,-13</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-9,9,-9</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-9,9,-9</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-5,9,-5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-5,9,-5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-41,9,-41</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-39,9,-39</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-39,9,-39</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-35,9,-35</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-35,9,-35</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-31,9,-31</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-31,9,-31</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-27,9,-27</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-27,9,-27</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-23,9,-23</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-23,9,-23</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-19,9,-19</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-19,9,-19</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-15,9,-15</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-15,9,-15</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-11,9,-11</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-11,9,-11</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-7,9,-7</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-7,9,-7</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>53.5,-36,53.5,-35.5</points>
<connection>
<GID>76</GID>
<name>clear</name></connection>
<connection>
<GID>145</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>54.5,-42,54.5,-42</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<connection>
<GID>144</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>52.5,-42,52.5,-42</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<connection>
<GID>145</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-9,251,53</points>
<intersection>-9 2</intersection>
<intersection>53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>251,53,258,53</points>
<connection>
<GID>85</GID>
<name>N_in0</name></connection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>250.5,-9,251,-9</points>
<connection>
<GID>147</GID>
<name>N_in1</name></connection>
<intersection>251 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251.5,-12,251.5,54</points>
<intersection>-12 2</intersection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>251.5,54,258,54</points>
<connection>
<GID>86</GID>
<name>N_in0</name></connection>
<intersection>251.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>250.5,-12,251.5,-12</points>
<connection>
<GID>148</GID>
<name>N_in1</name></connection>
<intersection>251.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>252.5,-15,252.5,55</points>
<intersection>-15 2</intersection>
<intersection>55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>252.5,55,258,55</points>
<connection>
<GID>87</GID>
<name>N_in0</name></connection>
<intersection>252.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>250.5,-15,252.5,-15</points>
<connection>
<GID>149</GID>
<name>N_in1</name></connection>
<intersection>252.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>253.5,-18,253.5,56</points>
<intersection>-18 2</intersection>
<intersection>56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>253.5,56,258,56</points>
<connection>
<GID>88</GID>
<name>N_in0</name></connection>
<intersection>253.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>250.5,-18,253.5,-18</points>
<connection>
<GID>150</GID>
<name>N_in1</name></connection>
<intersection>253.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-15,292,-15</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-13,286,-13</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-20,286,-17</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<connection>
<GID>162</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-16,286,-15</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<connection>
<GID>162</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-53,291,-51</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-51,291,-51</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-55,291,-55</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<connection>
<GID>176</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-59,290,-57</points>
<connection>
<GID>177</GID>
<name>OUT</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-57,291,-57</points>
<connection>
<GID>175</GID>
<name>IN_2</name></connection>
<intersection>290 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-64,291,-59</points>
<connection>
<GID>175</GID>
<name>IN_3</name></connection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>290,-64,291,-64</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-64,284,-64</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>297.5,8,297.5,8</points>
<connection>
<GID>193</GID>
<name>OUT</name></connection>
<connection>
<GID>194</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,1,290.5,5</points>
<connection>
<GID>193</GID>
<name>IN_3</name></connection>
<intersection>1 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>290,1,290.5,1</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,5,290,7</points>
<connection>
<GID>191</GID>
<name>OUT</name></connection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,7,290.5,7</points>
<connection>
<GID>193</GID>
<name>IN_2</name></connection>
<intersection>290 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268,-24,268,11</points>
<intersection>-24 2</intersection>
<intersection>-4 6</intersection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268,11,290.5,11</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>268 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>262,-24,291,-24</points>
<connection>
<GID>205</GID>
<name>N_in1</name></connection>
<intersection>268 0</intersection>
<intersection>291 21</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>268,-4,285.5,-4</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>268 0</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>291,-25,291,-24</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>-24 2</intersection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,4,284,4</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>284,0,284,0</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>267.5,-30,280,-30</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>267.5 50</intersection>
<intersection>280 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>280,-66,280,8</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>-66 47</intersection>
<intersection>-52 40</intersection>
<intersection>-48 22</intersection>
<intersection>-38 18</intersection>
<intersection>-30 1</intersection>
<intersection>-11 28</intersection>
<intersection>-7 38</intersection>
<intersection>8 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>280,8,284,8</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>280 5</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>280,-38,284,-38</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>280 5</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>280,-48,284,-48</points>
<connection>
<GID>173</GID>
<name>IN_2</name></connection>
<intersection>280 5</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>279.5,-11,280,-11</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>280 5</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>279.5,-7,280,-7</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>280 5</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>280,-52,284,-52</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>280 5</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>280,-66,284,-66</points>
<connection>
<GID>166</GID>
<name>IN_2</name></connection>
<intersection>280 5</intersection></hsegment>
<vsegment>
<ID>50</ID>
<points>267.5,-30,267.5,-27</points>
<intersection>-30 1</intersection>
<intersection>-27 51</intersection></vsegment>
<hsegment>
<ID>51</ID>
<points>262,-27,267.5,-27</points>
<connection>
<GID>202</GID>
<name>N_in1</name></connection>
<intersection>267.5 50</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-62,271,6</points>
<intersection>-62 41</intersection>
<intersection>-54 37</intersection>
<intersection>-50 35</intersection>
<intersection>-46 17</intersection>
<intersection>-36 30</intersection>
<intersection>-32 15</intersection>
<intersection>-25 45</intersection>
<intersection>-24 5</intersection>
<intersection>-13 39</intersection>
<intersection>-9 25</intersection>
<intersection>-5 11</intersection>
<intersection>2 1</intersection>
<intersection>6 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271,2,284,2</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>271,6,284,6</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>271,-24,280,-24</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>271,-5,279.5,-5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>271,-32,284,-32</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>271,-46,284,-46</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>271,-9,279.5,-9</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>271,-36,284,-36</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>271,-50,284,-50</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>271,-54,280,-54</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>271,-13,282,-13</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>271,-62,284,-62</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>262,-25,271,-25</points>
<connection>
<GID>204</GID>
<name>N_in1</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-64,276,10</points>
<intersection>-64 33</intersection>
<intersection>-58 28</intersection>
<intersection>-56 18</intersection>
<intersection>-44 16</intersection>
<intersection>-40 25</intersection>
<intersection>-34 12</intersection>
<intersection>-26 8</intersection>
<intersection>-19 26</intersection>
<intersection>-15 31</intersection>
<intersection>-2 1</intersection>
<intersection>4 2</intersection>
<intersection>10 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266.5,-2,285.5,-2</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>266.5 36</intersection>
<intersection>276 0</intersection>
<intersection>284 38</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,4,280,4</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>276,10,284,10</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>262,-26,284,-26</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<connection>
<GID>203</GID>
<name>N_in1</name></connection>
<intersection>266.5 36</intersection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>276,-34,280,-34</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>276,-44,280,-44</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>276,-56,284,-56</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>276,-40,284,-40</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>276,-19,280,-19</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>276,-58,284,-58</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>276,-15,280,-15</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>276,-64,280,-64</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>266.5,-26,266.5,-2</points>
<intersection>-26 8</intersection>
<intersection>-2 1</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>284,-28,284,-2</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>-2 1</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,9,290.5,9</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<connection>
<GID>197</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-27,290,-25</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>290,-27,291,-27</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>290 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-29,291,-29</points>
<connection>
<GID>199</GID>
<name>IN_2</name></connection>
<connection>
<GID>201</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-33,290.5,-31</points>
<intersection>-33 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-33,290.5,-33</points>
<connection>
<GID>184</GID>
<name>OUT</name></connection>
<intersection>290.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290.5,-31,291,-31</points>
<connection>
<GID>199</GID>
<name>IN_3</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-24,284,-24</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<connection>
<GID>200</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-30,284,-30</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<connection>
<GID>201</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-34,284,-34</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<connection>
<GID>184</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-28,298,-28</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<connection>
<GID>199</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296,-38,296,-38</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<connection>
<GID>188</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-41,290,-39</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<connection>
<GID>169</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-37,290,-37</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<connection>
<GID>171</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-42,284,-42</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-46,290,-46</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<connection>
<GID>190</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-44,284,-44</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-56,298,-56</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<connection>
<GID>189</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-54,284,-54</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-60,284,-60</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-5,292.5,-5</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<connection>
<GID>185</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-6,285.5,-6</points>
<connection>
<GID>180</GID>
<name>IN_2</name></connection>
<connection>
<GID>181</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-10,285.5,-8</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<connection>
<GID>180</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-97.5,292.5,-97.5</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<connection>
<GID>231</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,-95.5,286.5,-95.5</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,-102.5,286.5,-99.5</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<connection>
<GID>207</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,-98.5,286.5,-97.5</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<connection>
<GID>207</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-135.5,291.5,-133.5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>-133.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,-133.5,291.5,-133.5</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,-137.5,291.5,-137.5</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<connection>
<GID>221</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-141.5,290.5,-139.5</points>
<connection>
<GID>222</GID>
<name>OUT</name></connection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,-139.5,291.5,-139.5</points>
<connection>
<GID>220</GID>
<name>IN_2</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-146.5,291.5,-141.5</points>
<connection>
<GID>220</GID>
<name>IN_3</name></connection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>290.5,-146.5,291.5,-146.5</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-146.5,284.5,-146.5</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298,-74.5,298,-74.5</points>
<connection>
<GID>238</GID>
<name>OUT</name></connection>
<connection>
<GID>239</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-81.5,291,-77.5</points>
<connection>
<GID>238</GID>
<name>IN_3</name></connection>
<intersection>-81.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>290.5,-81.5,291,-81.5</points>
<connection>
<GID>237</GID>
<name>OUT</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-77.5,290.5,-75.5</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,-75.5,291,-75.5</points>
<connection>
<GID>238</GID>
<name>IN_2</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268.5,-106.5,268.5,-71.5</points>
<intersection>-106.5 2</intersection>
<intersection>-86.5 6</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,-71.5,291,-71.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>268.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>262.5,-106.5,291.5,-106.5</points>
<connection>
<GID>250</GID>
<name>N_in1</name></connection>
<intersection>268.5 0</intersection>
<intersection>291.5 21</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>268.5,-86.5,286,-86.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>268.5 0</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>291.5,-107.5,291.5,-106.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>-106.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-78.5,284.5,-78.5</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>284.5,-82.5,284.5,-82.5</points>
<connection>
<GID>237</GID>
<name>IN_1</name></connection>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>268,-112.5,280.5,-112.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>268 50</intersection>
<intersection>280.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>280.5,-148.5,280.5,-74.5</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>-148.5 47</intersection>
<intersection>-134.5 40</intersection>
<intersection>-130.5 22</intersection>
<intersection>-120.5 18</intersection>
<intersection>-112.5 1</intersection>
<intersection>-93.5 28</intersection>
<intersection>-89.5 38</intersection>
<intersection>-74.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>280.5,-74.5,284.5,-74.5</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>280.5 5</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>280.5,-120.5,284.5,-120.5</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>280.5 5</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>280.5,-130.5,284.5,-130.5</points>
<connection>
<GID>218</GID>
<name>IN_2</name></connection>
<intersection>280.5 5</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>280,-93.5,280.5,-93.5</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<intersection>280.5 5</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>280,-89.5,280.5,-89.5</points>
<connection>
<GID>226</GID>
<name>IN_1</name></connection>
<intersection>280.5 5</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>280.5,-134.5,284.5,-134.5</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>280.5 5</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>280.5,-148.5,284.5,-148.5</points>
<connection>
<GID>211</GID>
<name>IN_2</name></connection>
<intersection>280.5 5</intersection></hsegment>
<vsegment>
<ID>50</ID>
<points>268,-112.5,268,-109.5</points>
<intersection>-112.5 1</intersection>
<intersection>-109.5 51</intersection></vsegment>
<hsegment>
<ID>51</ID>
<points>262.5,-109.5,268,-109.5</points>
<connection>
<GID>247</GID>
<name>N_in1</name></connection>
<intersection>268 50</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-144.5,271.5,-76.5</points>
<intersection>-144.5 41</intersection>
<intersection>-136.5 37</intersection>
<intersection>-132.5 35</intersection>
<intersection>-128.5 17</intersection>
<intersection>-118.5 30</intersection>
<intersection>-114.5 15</intersection>
<intersection>-107.5 45</intersection>
<intersection>-106.5 5</intersection>
<intersection>-95.5 39</intersection>
<intersection>-91.5 25</intersection>
<intersection>-87.5 11</intersection>
<intersection>-80.5 1</intersection>
<intersection>-76.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271.5,-80.5,284.5,-80.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>271.5,-76.5,284.5,-76.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>271.5,-106.5,280.5,-106.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>271.5,-87.5,280,-87.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>271.5,-114.5,284.5,-114.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>271.5,-128.5,284.5,-128.5</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>271.5,-91.5,280,-91.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>271.5,-118.5,284.5,-118.5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>271.5,-132.5,284.5,-132.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>271.5,-136.5,280.5,-136.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>271.5,-95.5,282.5,-95.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>271.5,-144.5,284.5,-144.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>262.5,-107.5,271.5,-107.5</points>
<connection>
<GID>249</GID>
<name>N_in1</name></connection>
<intersection>271.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276.5,-146.5,276.5,-72.5</points>
<intersection>-146.5 33</intersection>
<intersection>-140.5 28</intersection>
<intersection>-138.5 18</intersection>
<intersection>-126.5 16</intersection>
<intersection>-122.5 25</intersection>
<intersection>-116.5 12</intersection>
<intersection>-108.5 8</intersection>
<intersection>-101.5 26</intersection>
<intersection>-97.5 31</intersection>
<intersection>-84.5 1</intersection>
<intersection>-78.5 2</intersection>
<intersection>-72.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267,-84.5,286,-84.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>267 36</intersection>
<intersection>276.5 0</intersection>
<intersection>284.5 38</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276.5,-78.5,280.5,-78.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>276.5,-72.5,284.5,-72.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>262.5,-108.5,284.5,-108.5</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<connection>
<GID>248</GID>
<name>N_in1</name></connection>
<intersection>267 36</intersection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>276.5,-116.5,280.5,-116.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>276.5,-126.5,280.5,-126.5</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>276.5,-138.5,284.5,-138.5</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>276.5,-122.5,284.5,-122.5</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>276.5,-101.5,280.5,-101.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>276.5,-140.5,284.5,-140.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>276.5,-97.5,280.5,-97.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>276.5,-146.5,280.5,-146.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>267,-108.5,267,-84.5</points>
<intersection>-108.5 8</intersection>
<intersection>-84.5 1</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>284.5,-110.5,284.5,-84.5</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>-84.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,-73.5,291,-73.5</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<connection>
<GID>242</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-109.5,290.5,-107.5</points>
<connection>
<GID>245</GID>
<name>OUT</name></connection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>290.5,-109.5,291.5,-109.5</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,-111.5,291.5,-111.5</points>
<connection>
<GID>244</GID>
<name>IN_2</name></connection>
<connection>
<GID>246</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-115.5,291,-113.5</points>
<intersection>-115.5 1</intersection>
<intersection>-113.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,-115.5,291,-115.5</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291,-113.5,291.5,-113.5</points>
<connection>
<GID>244</GID>
<name>IN_3</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-106.5,284.5,-106.5</points>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection>
<connection>
<GID>245</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-112.5,284.5,-112.5</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<connection>
<GID>246</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-116.5,284.5,-116.5</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<connection>
<GID>229</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-110.5,298.5,-110.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<connection>
<GID>244</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,-120.5,296.5,-120.5</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<connection>
<GID>233</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-123.5,290.5,-121.5</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<connection>
<GID>214</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-119.5,290.5,-119.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<connection>
<GID>216</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-124.5,284.5,-124.5</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-128.5,290.5,-128.5</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<connection>
<GID>235</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-126.5,284.5,-126.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298.5,-138.5,298.5,-138.5</points>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<connection>
<GID>234</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-136.5,284.5,-136.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-142.5,284.5,-142.5</points>
<connection>
<GID>222</GID>
<name>IN_1</name></connection>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>293,-87.5,293.5,-87.5</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<connection>
<GID>230</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-88.5,286,-88.5</points>
<connection>
<GID>225</GID>
<name>IN_2</name></connection>
<connection>
<GID>226</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-92.5,286,-90.5</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<connection>
<GID>225</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255,-27,255,-23</points>
<intersection>-27 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-23,255,-23</points>
<connection>
<GID>151</GID>
<name>N_in1</name></connection>
<intersection>255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>255,-27,260,-27</points>
<connection>
<GID>202</GID>
<name>N_in0</name></connection>
<intersection>255 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>250.5,-26,260,-26</points>
<connection>
<GID>152</GID>
<name>N_in1</name></connection>
<connection>
<GID>203</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255,-29,255,-25</points>
<intersection>-29 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-29,255,-29</points>
<connection>
<GID>153</GID>
<name>N_in1</name></connection>
<intersection>255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>255,-25,260,-25</points>
<connection>
<GID>204</GID>
<name>N_in0</name></connection>
<intersection>255 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255,-32,255,-24</points>
<intersection>-32 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-32,255,-32</points>
<connection>
<GID>154</GID>
<name>N_in1</name></connection>
<intersection>255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>255,-24,260,-24</points>
<connection>
<GID>205</GID>
<name>N_in0</name></connection>
<intersection>255 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255.5,-109.5,255.5,-36</points>
<intersection>-109.5 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-36,255.5,-36</points>
<connection>
<GID>155</GID>
<name>N_in1</name></connection>
<intersection>255.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>255.5,-109.5,260.5,-109.5</points>
<connection>
<GID>247</GID>
<name>N_in0</name></connection>
<intersection>255.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255.5,-108.5,255.5,-39</points>
<intersection>-108.5 1</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-108.5,260.5,-108.5</points>
<connection>
<GID>248</GID>
<name>N_in0</name></connection>
<intersection>255.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>250.5,-39,255.5,-39</points>
<connection>
<GID>156</GID>
<name>N_in1</name></connection>
<intersection>255.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255.5,-107.5,255.5,-42</points>
<intersection>-107.5 2</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-42,255.5,-42</points>
<connection>
<GID>157</GID>
<name>N_in1</name></connection>
<intersection>255.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>255.5,-107.5,260.5,-107.5</points>
<connection>
<GID>249</GID>
<name>N_in0</name></connection>
<intersection>255.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255.5,-106.5,255.5,-45</points>
<intersection>-106.5 1</intersection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-106.5,260.5,-106.5</points>
<connection>
<GID>250</GID>
<name>N_in0</name></connection>
<intersection>255.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>250.5,-45,255.5,-45</points>
<connection>
<GID>158</GID>
<name>N_in1</name></connection>
<intersection>255.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-18,242,-9</points>
<intersection>-18 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242,-9,248.5,-9</points>
<connection>
<GID>147</GID>
<name>N_in0</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235.5,-18,242,-18</points>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-16,242,-12</points>
<intersection>-16 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242,-12,248.5,-12</points>
<connection>
<GID>148</GID>
<name>N_in0</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235.5,-16,242,-16</points>
<connection>
<GID>160</GID>
<name>OUT_1</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-15,242,-14</points>
<intersection>-15 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242,-15,248.5,-15</points>
<connection>
<GID>149</GID>
<name>N_in0</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235.5,-14,242,-14</points>
<connection>
<GID>160</GID>
<name>OUT_2</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-18,242,-12</points>
<intersection>-18 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242,-18,248.5,-18</points>
<connection>
<GID>150</GID>
<name>N_in0</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235.5,-12,242,-12</points>
<connection>
<GID>160</GID>
<name>OUT_3</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,46.3715,715.223,-326.526</PageViewport></page 2>
<page 3>
<PageViewport>0,46.3715,715.223,-326.526</PageViewport></page 3>
<page 4>
<PageViewport>0,46.3715,715.223,-326.526</PageViewport></page 4>
<page 5>
<PageViewport>0,46.3715,715.223,-326.526</PageViewport></page 5>
<page 6>
<PageViewport>0,46.3715,715.223,-326.526</PageViewport></page 6>
<page 7>
<PageViewport>0,46.3715,715.223,-326.526</PageViewport></page 7>
<page 8>
<PageViewport>0,46.3715,715.223,-326.526</PageViewport></page 8>
<page 9>
<PageViewport>0,46.3715,715.223,-326.526</PageViewport></page 9></circuit>