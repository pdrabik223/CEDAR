<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-0.199999,-0.1,177.6,-92.8</PageViewport>
<gate>
<ID>2</ID>
<type>DD_KEYPAD_HEX</type>
<position>5.5,-13</position>
<output>
<ID>OUT_0</ID>30 </output>
<output>
<ID>OUT_1</ID>32 </output>
<output>
<ID>OUT_2</ID>33 </output>
<output>
<ID>OUT_3</ID>34 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>4</ID>
<type>DD_KEYPAD_HEX</type>
<position>5.5,-25.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<output>
<ID>OUT_1</ID>42 </output>
<output>
<ID>OUT_2</ID>47 </output>
<output>
<ID>OUT_3</ID>56 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>6</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>125.5,-22.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_2</ID>52 </input>
<input>
<ID>IN_3</ID>77 </input>
<input>
<ID>IN_4</ID>78 </input>
<input>
<ID>IN_5</ID>79 </input>
<input>
<ID>IN_6</ID>80 </input>
<input>
<ID>IN_7</ID>84 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 16</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>20.5,-20.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>6,-4</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>5,-33.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_AND2</type>
<position>19,-14.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND2</type>
<position>19,-10.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND2</type>
<position>19,-6.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_FULLADDER_4BIT</type>
<position>41.5,-10.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>41 </input>
<input>
<ID>IN_B_1</ID>37 </input>
<input>
<ID>IN_B_2</ID>36 </input>
<input>
<ID>IN_B_3</ID>35 </input>
<output>
<ID>OUT_0</ID>46 </output>
<output>
<ID>OUT_1</ID>45 </output>
<output>
<ID>OUT_2</ID>44 </output>
<output>
<ID>OUT_3</ID>43 </output>
<output>
<ID>overflow</ID>83 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_AND2</type>
<position>30.5,-31.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>30.5,-35.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>30.5,-39.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_AND2</type>
<position>30.5,-43.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AE_FULLADDER_4BIT</type>
<position>58.5,-11</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>49 </input>
<input>
<ID>IN_2</ID>50 </input>
<input>
<ID>IN_3</ID>51 </input>
<input>
<ID>IN_B_1</ID>46 </input>
<input>
<ID>IN_B_2</ID>45 </input>
<input>
<ID>IN_B_3</ID>44 </input>
<output>
<ID>OUT_0</ID>55 </output>
<output>
<ID>OUT_1</ID>54 </output>
<output>
<ID>OUT_2</ID>53 </output>
<output>
<ID>OUT_3</ID>52 </output>
<input>
<ID>carry_in</ID>83 </input>
<output>
<ID>overflow</ID>82 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>55,-29</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>55,-33</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>55,-37</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>55,-41</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_FULLADDER_4BIT</type>
<position>71,-36</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>60 </input>
<input>
<ID>IN_B_1</ID>55 </input>
<input>
<ID>IN_B_2</ID>54 </input>
<input>
<ID>IN_B_3</ID>53 </input>
<output>
<ID>OUT_0</ID>80 </output>
<output>
<ID>OUT_1</ID>79 </output>
<output>
<ID>OUT_2</ID>78 </output>
<output>
<ID>OUT_3</ID>77 </output>
<input>
<ID>carry_in</ID>82 </input>
<output>
<ID>overflow</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_AND2</type>
<position>54.5,-48</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>54.5,-52</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND2</type>
<position>54.5,-56</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_AND2</type>
<position>54.5,-60</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>13</ID>
<points>14.5,-28.5,14.5,-7.5</points>
<intersection>-28.5 14</intersection>
<intersection>-21.5 21</intersection>
<intersection>-15.5 23</intersection>
<intersection>-11.5 25</intersection>
<intersection>-7.5 27</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>10.5,-28.5,14.5,-28.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>14.5 13</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>14.5,-21.5,17.5,-21.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>14.5 13</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>14.5,-15.5,16,-15.5</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>14.5 13</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>14.5,-11.5,16,-11.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>14.5 13</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>14.5,-7.5,16,-7.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>14.5 13</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>12.5,-19.5,17.5,-19.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>12.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>12.5,-59,12.5,-16</points>
<intersection>-59 14</intersection>
<intersection>-42.5 10</intersection>
<intersection>-19.5 2</intersection>
<intersection>-16 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>12.5,-42.5,52,-42.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>12.5 8</intersection>
<intersection>52 12</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>10.5,-16,12.5,-16</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>12.5 8</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>52,-42.5,52,-40</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-42.5 10</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>12.5,-59,51.5,-59</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>12.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>23.5,-25.5,120.5,-25.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>23.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23.5,-25.5,23.5,-20.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>-25.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10.5,-13.5,16,-13.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>10.5 9</intersection>
<intersection>13.5 10</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>10.5,-14,10.5,-13.5</points>
<intersection>-14 15</intersection>
<intersection>-13.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>13.5,-38.5,13.5,-13.5</points>
<intersection>-38.5 11</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>13.5,-38.5,52,-38.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>13.5 10</intersection>
<intersection>14 13</intersection>
<intersection>52 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>52,-38.5,52,-36</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-38.5 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>14,-55,14,-38.5</points>
<intersection>-55 14</intersection>
<intersection>-38.5 11</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>14,-55,51.5,-55</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>14 13</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>10.5,-14,10.5,-14</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>10.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-34.5,13,-9.5</points>
<intersection>-34.5 3</intersection>
<intersection>-12 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-12,13,-12</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-9.5,16,-9.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>13,-34.5,52,-34.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection>
<intersection>16.5 5</intersection>
<intersection>52 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>52,-34.5,52,-32</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-34.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>16.5,-51,16.5,-34.5</points>
<intersection>-51 6</intersection>
<intersection>-34.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>16.5,-51,51.5,-51</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>16.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-30.5,12.5,-5.5</points>
<intersection>-30.5 3</intersection>
<intersection>-10 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-10,12.5,-10</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-5.5,16,-5.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>12.5,-30.5,52,-30.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection>
<intersection>21 5</intersection>
<intersection>52 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>52,-30.5,52,-28</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>-30.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>21,-47,21,-30.5</points>
<intersection>-47 6</intersection>
<intersection>-30.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>21,-47,51.5,-47</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>21 5</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-14.5,23.5,-8.5</points>
<intersection>-14.5 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-8.5,37.5,-8.5</points>
<connection>
<GID>31</GID>
<name>IN_B_3</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-14.5,23.5,-14.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-7.5,37.5,-7.5</points>
<connection>
<GID>31</GID>
<name>IN_B_2</name></connection>
<intersection>22 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22,-10.5,22,-7.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>-7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-6.5,37.5,-6.5</points>
<connection>
<GID>31</GID>
<name>IN_B_1</name></connection>
<intersection>22 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>22,-6.5,22,-6.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>-6.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-31.5,35,-12.5</points>
<intersection>-31.5 2</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-12.5,37.5,-12.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-31.5,35,-31.5</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-35.5,36,-13.5</points>
<intersection>-35.5 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-13.5,37.5,-13.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-35.5,36,-35.5</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-39.5,37,-14.5</points>
<intersection>-39.5 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-39.5,37,-39.5</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-14.5,37.5,-14.5</points>
<connection>
<GID>31</GID>
<name>IN_2</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-43.5,37,-15.5</points>
<intersection>-43.5 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-43.5,37,-43.5</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-15.5,37.5,-15.5</points>
<connection>
<GID>31</GID>
<name>IN_3</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-44.5,19,-26.5</points>
<intersection>-44.5 8</intersection>
<intersection>-40.5 6</intersection>
<intersection>-36.5 4</intersection>
<intersection>-32.5 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-32.5,27.5,-32.5</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10.5,-26.5,19,-26.5</points>
<connection>
<GID>4</GID>
<name>OUT_1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>19,-36.5,27.5,-36.5</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>19,-40.5,27.5,-40.5</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>19,-44.5,27.5,-44.5</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-24.5,45.5,-12</points>
<connection>
<GID>31</GID>
<name>OUT_3</name></connection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-24.5,120.5,-24.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-11,50,-9</points>
<intersection>-11 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-9,54.5,-9</points>
<connection>
<GID>40</GID>
<name>IN_B_3</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-11,50,-11</points>
<connection>
<GID>31</GID>
<name>OUT_2</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-10,50,-8</points>
<intersection>-10 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-8,54.5,-8</points>
<connection>
<GID>40</GID>
<name>IN_B_2</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-10,50,-10</points>
<connection>
<GID>31</GID>
<name>OUT_1</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-9,50,-7</points>
<intersection>-9 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-7,54.5,-7</points>
<connection>
<GID>40</GID>
<name>IN_B_1</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-9,50,-9</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-42,43.5,-24.5</points>
<intersection>-42 8</intersection>
<intersection>-38 6</intersection>
<intersection>-34 4</intersection>
<intersection>-30 1</intersection>
<intersection>-24.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-30,52,-30</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>43.5,-34,52,-34</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>43.5,-38,52,-38</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>43.5,-42,52,-42</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>10.5,-24.5,43.5,-24.5</points>
<connection>
<GID>4</GID>
<name>OUT_2</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-29,56,-13</points>
<intersection>-29 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-13,56,-13</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-29,58,-29</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-33,56,-14</points>
<intersection>-33 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-14,56,-14</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-33,58,-33</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-37,56,-15</points>
<intersection>-37 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-15,56,-15</points>
<connection>
<GID>40</GID>
<name>IN_2</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-37,58,-37</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-41,56,-16</points>
<intersection>-41 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-16,56,-16</points>
<connection>
<GID>40</GID>
<name>IN_3</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-41,58,-41</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-23.5,65,-12.5</points>
<intersection>-23.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,-23.5,120.5,-23.5</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-12.5,65,-12.5</points>
<connection>
<GID>40</GID>
<name>OUT_3</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-34,64.5,-11.5</points>
<intersection>-34 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-11.5,64.5,-11.5</points>
<connection>
<GID>40</GID>
<name>OUT_2</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-34,67,-34</points>
<connection>
<GID>45</GID>
<name>IN_B_3</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-33,64.5,-10.5</points>
<intersection>-33 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-10.5,64.5,-10.5</points>
<connection>
<GID>40</GID>
<name>OUT_1</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-33,67,-33</points>
<connection>
<GID>45</GID>
<name>IN_B_2</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-32,64.5,-9.5</points>
<intersection>-32 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-9.5,64.5,-9.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-32,67,-32</points>
<connection>
<GID>45</GID>
<name>IN_B_1</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-61,11.5,-22.5</points>
<intersection>-61 13</intersection>
<intersection>-57 14</intersection>
<intersection>-53 15</intersection>
<intersection>-49 16</intersection>
<intersection>-22.5 17</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>11.5,-61,51.5,-61</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>11.5,-57,51.5,-57</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>11.5,-53,51.5,-53</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>11.5,-49,51.5,-49</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>10.5,-22.5,11.5,-22.5</points>
<connection>
<GID>4</GID>
<name>OUT_3</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-48,61.5,-38</points>
<intersection>-48 2</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-38,67,-38</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-48,61.5,-48</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-52,62,-39</points>
<intersection>-52 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-39,67,-39</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-52,62,-52</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-56,62,-40</points>
<intersection>-56 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-40,67,-40</points>
<connection>
<GID>45</GID>
<name>IN_2</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-56,62,-56</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-60,62,-41</points>
<intersection>-60 2</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-41,67,-41</points>
<connection>
<GID>45</GID>
<name>IN_3</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-60,62,-60</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-37.5,79,-22.5</points>
<intersection>-37.5 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-22.5,120.5,-22.5</points>
<connection>
<GID>6</GID>
<name>IN_3</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-37.5,79,-37.5</points>
<connection>
<GID>45</GID>
<name>OUT_3</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-36.5,77.5,-21.5</points>
<intersection>-36.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-21.5,120.5,-21.5</points>
<connection>
<GID>6</GID>
<name>IN_4</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-36.5,77.5,-36.5</points>
<connection>
<GID>45</GID>
<name>OUT_2</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-35.5,76.5,-20.5</points>
<intersection>-35.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-20.5,120.5,-20.5</points>
<connection>
<GID>6</GID>
<name>IN_5</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-35.5,76.5,-35.5</points>
<connection>
<GID>45</GID>
<name>OUT_1</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-34.5,75.5,-19.5</points>
<intersection>-34.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-19.5,120.5,-19.5</points>
<connection>
<GID>6</GID>
<name>IN_6</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-34.5,75.5,-34.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-23.5,59.5,-19</points>
<connection>
<GID>40</GID>
<name>overflow</name></connection>
<intersection>-23.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>70,-28,70,-23.5</points>
<connection>
<GID>45</GID>
<name>carry_in</name></connection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59.5,-23.5,70,-23.5</points>
<intersection>59.5 0</intersection>
<intersection>70 1</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-10.5,57.5,-3</points>
<connection>
<GID>40</GID>
<name>carry_in</name></connection>
<intersection>-10.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>42.5,-18.5,42.5,-10.5</points>
<connection>
<GID>31</GID>
<name>overflow</name></connection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-10.5,57.5,-10.5</points>
<intersection>42.5 1</intersection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-44,83.5,-18.5</points>
<intersection>-44 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-18.5,120.5,-18.5</points>
<connection>
<GID>6</GID>
<name>IN_7</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-44,83.5,-44</points>
<connection>
<GID>45</GID>
<name>overflow</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 9></circuit>