<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-76.8872,115.987,211.145,-34.1852</PageViewport>
<gate>
<ID>593</ID>
<type>GA_LED</type>
<position>2,71</position>
<input>
<ID>N_in0</ID>366 </input>
<gparam>LED_BOX -30,-20,30,20</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>594</ID>
<type>AA_TOGGLE</type>
<position>-32.5,71</position>
<output>
<ID>OUT_0</ID>366 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>CC_PULSE</type>
<position>-3.5,17</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>27</ID>
<type>CC_PULSE</type>
<position>0.5,39.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>28</ID>
<type>CC_PULSE</type>
<position>-3.5,39.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>29</ID>
<type>CC_PULSE</type>
<position>-7.5,39.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>30</ID>
<type>CC_PULSE</type>
<position>0.5,32</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>31</ID>
<type>CC_PULSE</type>
<position>-3.5,32</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>32</ID>
<type>CC_PULSE</type>
<position>-7.5,32</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>33</ID>
<type>CC_PULSE</type>
<position>0.5,24.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>34</ID>
<type>CC_PULSE</type>
<position>-3.5,24.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>35</ID>
<type>CC_PULSE</type>
<position>-7.5,24.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>-7.5,43.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>616</ID>
<type>GA_LED</type>
<position>21.5,79</position>
<input>
<ID>N_in2</ID>370 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>-3.5,43.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>617</ID>
<type>GA_LED</type>
<position>15,72.5</position>
<input>
<ID>N_in0</ID>371 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>0.5,43.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>618</ID>
<type>GA_LED</type>
<position>8.5,79</position>
<input>
<ID>N_in2</ID>367 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>-7.5,36</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>619</ID>
<type>GA_LED</type>
<position>15,85.5</position>
<input>
<ID>N_in2</ID>368 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>-3.5,36</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>620</ID>
<type>GA_LED</type>
<position>21.5,66</position>
<input>
<ID>N_in3</ID>373 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>41</ID>
<type>DE_TO</type>
<position>0.5,36</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>621</ID>
<type>GA_LED</type>
<position>8.5,66</position>
<input>
<ID>N_in0</ID>372 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>-7.5,28.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>622</ID>
<type>GA_LED</type>
<position>15,59.5</position>
<input>
<ID>N_in2</ID>374 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>-3.5,28.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>0.5,28.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>-3.5,21</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>644</ID>
<type>GA_LED</type>
<position>4,79</position>
<input>
<ID>N_in2</ID>377 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>645</ID>
<type>GA_LED</type>
<position>-2.5,72.5</position>
<input>
<ID>N_in0</ID>378 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>646</ID>
<type>GA_LED</type>
<position>-9,79</position>
<input>
<ID>N_in2</ID>375 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>647</ID>
<type>GA_LED</type>
<position>-2.5,85.5</position>
<input>
<ID>N_in2</ID>376 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>648</ID>
<type>GA_LED</type>
<position>4,66</position>
<input>
<ID>N_in3</ID>380 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>649</ID>
<type>GA_LED</type>
<position>-9,66</position>
<input>
<ID>N_in0</ID>379 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>650</ID>
<type>GA_LED</type>
<position>-2.5,59.5</position>
<input>
<ID>N_in2</ID>381 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>651</ID>
<type>DA_FROM</type>
<position>-8,97</position>
<input>
<ID>IN_0</ID>381 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b7</lparam></gate>
<gate>
<ID>652</ID>
<type>DA_FROM</type>
<position>-6,97</position>
<input>
<ID>IN_0</ID>380 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b6</lparam></gate>
<gate>
<ID>653</ID>
<type>DA_FROM</type>
<position>-4,97</position>
<input>
<ID>IN_0</ID>379 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b5</lparam></gate>
<gate>
<ID>654</ID>
<type>DA_FROM</type>
<position>-2,97</position>
<input>
<ID>IN_0</ID>378 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b4</lparam></gate>
<gate>
<ID>655</ID>
<type>DA_FROM</type>
<position>0,97</position>
<input>
<ID>IN_0</ID>377 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b3</lparam></gate>
<gate>
<ID>656</ID>
<type>DA_FROM</type>
<position>2,97</position>
<input>
<ID>IN_0</ID>376 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b2</lparam></gate>
<gate>
<ID>77</ID>
<type>CC_PULSE</type>
<position>10,17</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>657</ID>
<type>DA_FROM</type>
<position>4,97</position>
<input>
<ID>IN_0</ID>375 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID b1</lparam></gate>
<gate>
<ID>78</ID>
<type>DE_TO</type>
<position>10,21</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>658</ID>
<type>GA_LED</type>
<position>-13,79</position>
<input>
<ID>N_in2</ID>384 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>659</ID>
<type>GA_LED</type>
<position>-19.5,72.5</position>
<input>
<ID>N_in0</ID>385 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>660</ID>
<type>GA_LED</type>
<position>-26,79</position>
<input>
<ID>N_in2</ID>382 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>661</ID>
<type>GA_LED</type>
<position>-19.5,85.5</position>
<input>
<ID>N_in2</ID>383 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>662</ID>
<type>GA_LED</type>
<position>-13,66</position>
<input>
<ID>N_in3</ID>387 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>663</ID>
<type>GA_LED</type>
<position>-26,66</position>
<input>
<ID>N_in0</ID>386 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>664</ID>
<type>GA_LED</type>
<position>-19.5,59.5</position>
<input>
<ID>N_in2</ID>388 </input>
<gparam>LED_BOX -5.4,-1.1,5.4,1.1</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>665</ID>
<type>DA_FROM</type>
<position>-25,97</position>
<input>
<ID>IN_0</ID>388 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c7</lparam></gate>
<gate>
<ID>666</ID>
<type>DA_FROM</type>
<position>-23,97</position>
<input>
<ID>IN_0</ID>387 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c6</lparam></gate>
<gate>
<ID>667</ID>
<type>DA_FROM</type>
<position>-21,97</position>
<input>
<ID>IN_0</ID>386 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c5</lparam></gate>
<gate>
<ID>668</ID>
<type>DA_FROM</type>
<position>-19,97</position>
<input>
<ID>IN_0</ID>385 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c4</lparam></gate>
<gate>
<ID>669</ID>
<type>DA_FROM</type>
<position>-17,97</position>
<input>
<ID>IN_0</ID>384 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c3</lparam></gate>
<gate>
<ID>670</ID>
<type>DA_FROM</type>
<position>-15,97</position>
<input>
<ID>IN_0</ID>383 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c2</lparam></gate>
<gate>
<ID>671</ID>
<type>DA_FROM</type>
<position>-13,97</position>
<input>
<ID>IN_0</ID>382 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID c1</lparam></gate>
<gate>
<ID>561</ID>
<type>DA_FROM</type>
<position>9.5,97</position>
<input>
<ID>IN_0</ID>374 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a7</lparam></gate>
<gate>
<ID>562</ID>
<type>DA_FROM</type>
<position>11.5,97</position>
<input>
<ID>IN_0</ID>373 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a6</lparam></gate>
<gate>
<ID>563</ID>
<type>DA_FROM</type>
<position>13.5,97</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a5</lparam></gate>
<gate>
<ID>564</ID>
<type>DA_FROM</type>
<position>15.5,97</position>
<input>
<ID>IN_0</ID>371 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a4</lparam></gate>
<gate>
<ID>571</ID>
<type>DA_FROM</type>
<position>17.5,97</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a3</lparam></gate>
<gate>
<ID>572</ID>
<type>DA_FROM</type>
<position>19.5,97</position>
<input>
<ID>IN_0</ID>368 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a2</lparam></gate>
<gate>
<ID>573</ID>
<type>DA_FROM</type>
<position>21.5,97</position>
<input>
<ID>IN_0</ID>367 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a1</lparam></gate>
<wire>
<ID>386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,65,-25,73.5</points>
<intersection>65 4</intersection>
<intersection>73.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-14,73.5,-14,95</points>
<intersection>73.5 2</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-25,73.5,-14,73.5</points>
<intersection>-25 0</intersection>
<intersection>-14 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-21,95,-14,95</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-26,65,-25,65</points>
<connection>
<GID>663</GID>
<name>N_in0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,66,-14,95</points>
<connection>
<GID>662</GID>
<name>N_in3</name></connection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-23,95,-14,95</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,60.5,-14,95</points>
<intersection>60.5 4</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-25,95,-14,95</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-19.5,60.5,-14,60.5</points>
<connection>
<GID>664</GID>
<name>N_in2</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,41.5,-7.5,41.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,41.5,-3.5,41.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,41.5,0.5,41.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,34,-7.5,34</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,34,-3.5,34</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>0.5,34,0.5,34</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<connection>
<GID>41</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,26.5,-7.5,26.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,26.5,-3.5,26.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,26.5,0.5,26.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<connection>
<GID>44</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,19,-3.5,19</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,19,10,19</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-30.5,71,1,71</points>
<connection>
<GID>594</GID>
<name>OUT_0</name></connection>
<connection>
<GID>593</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,73.5,20.5,95</points>
<intersection>73.5 1</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,73.5,20.5,73.5</points>
<intersection>9.5 2</intersection>
<intersection>20.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>9.5,73.5,9.5,79</points>
<connection>
<GID>618</GID>
<name>N_in2</name></connection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>20.5,95,21.5,95</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,86.5,20.5,95</points>
<intersection>86.5 3</intersection>
<intersection>95 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>15,86.5,20.5,86.5</points>
<connection>
<GID>619</GID>
<name>N_in2</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>19.5,95,20.5,95</points>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,79,20.5,95</points>
<intersection>79 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,79,22.5,79</points>
<connection>
<GID>616</GID>
<name>N_in2</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,95,20.5,95</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,72.5,20.5,95</points>
<intersection>72.5 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,72.5,20.5,72.5</points>
<connection>
<GID>617</GID>
<name>N_in0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,95,20.5,95</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,65,9.5,71.5</points>
<intersection>65 4</intersection>
<intersection>71.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>20.5,71.5,20.5,95</points>
<intersection>71.5 2</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9.5,71.5,20.5,71.5</points>
<intersection>9.5 0</intersection>
<intersection>20.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>13.5,95,20.5,95</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<intersection>20.5 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>8.5,65,9.5,65</points>
<connection>
<GID>621</GID>
<name>N_in0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,66,20.5,95</points>
<connection>
<GID>620</GID>
<name>N_in3</name></connection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11.5,95,20.5,95</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,60.5,20.5,95</points>
<intersection>60.5 4</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>9.5,95,20.5,95</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>15,60.5,20.5,60.5</points>
<connection>
<GID>622</GID>
<name>N_in2</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,73.5,3,95</points>
<intersection>73.5 1</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,73.5,3,73.5</points>
<intersection>-8 2</intersection>
<intersection>3 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-8,73.5,-8,79</points>
<connection>
<GID>646</GID>
<name>N_in2</name></connection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>3,95,4,95</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,86.5,3,95</points>
<intersection>86.5 3</intersection>
<intersection>95 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2.5,86.5,3,86.5</points>
<connection>
<GID>647</GID>
<name>N_in2</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>2,95,3,95</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,79,3,95</points>
<intersection>79 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,79,5,79</points>
<connection>
<GID>644</GID>
<name>N_in2</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.30078e-008,95,3,95</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,72.5,3,95</points>
<intersection>72.5 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,72.5,3,72.5</points>
<connection>
<GID>645</GID>
<name>N_in0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,95,3,95</points>
<connection>
<GID>654</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,65,-8,73.5</points>
<intersection>65 4</intersection>
<intersection>73.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>3,73.5,3,95</points>
<intersection>73.5 2</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8,73.5,3,73.5</points>
<intersection>-8 0</intersection>
<intersection>3 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4,95,3,95</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>3 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-9,65,-8,65</points>
<connection>
<GID>649</GID>
<name>N_in0</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,66,3,95</points>
<connection>
<GID>648</GID>
<name>N_in3</name></connection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-6,95,3,95</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,60.5,3,95</points>
<intersection>60.5 4</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-8,95,3,95</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-2.5,60.5,3,60.5</points>
<connection>
<GID>650</GID>
<name>N_in2</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,73.5,-14,95</points>
<intersection>73.5 1</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,73.5,-14,73.5</points>
<intersection>-25 2</intersection>
<intersection>-14 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-25,73.5,-25,79</points>
<connection>
<GID>660</GID>
<name>N_in2</name></connection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-14,95,-13,95</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,86.5,-14,95</points>
<intersection>86.5 3</intersection>
<intersection>95 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,86.5,-14,86.5</points>
<connection>
<GID>661</GID>
<name>N_in2</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-15,95,-14,95</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,79,-14,95</points>
<intersection>79 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,79,-12,79</points>
<connection>
<GID>658</GID>
<name>N_in2</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-17,95,-14,95</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,72.5,-14,95</points>
<intersection>72.5 1</intersection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-18.5,72.5,-14,72.5</points>
<connection>
<GID>659</GID>
<name>N_in0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19,95,-14,95</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-24.0855,59.77,331.916,-125.839</PageViewport>
<gate>
<ID>1</ID>
<type>BM_NORX2</type>
<position>231,30</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_OR3</type>
<position>233,66</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>3 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_SMALL_INVERTER</type>
<position>228,68</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>BM_NORX2</type>
<position>227,65</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,57</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND3</type>
<position>231,17</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>26 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,51</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,47</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_OR2</type>
<position>237,43</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>231,40</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>BM_NORX2</type>
<position>231,44</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,39</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_OR3</type>
<position>231,35</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>27 </input>
<input>
<ID>IN_2</ID>26 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,37</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>15</ID>
<type>AE_OR4</type>
<position>238,25</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>231,26</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_AND2</type>
<position>231,22</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,27</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,21</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_OR4</type>
<position>232.5,76</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>23 </input>
<input>
<ID>IN_2</ID>71 </input>
<input>
<ID>IN_3</ID>72 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>21</ID>
<type>BM_NORX2</type>
<position>226.5,75</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>226.5,71</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,17</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>231,48</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>DE_TO</type>
<position>238.5,76</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a2</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>238,66</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a3</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>244,53</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a4</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>242,43</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a5</lparam></gate>
<gate>
<ID>49</ID>
<type>DE_TO</type>
<position>244,25</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a7</lparam></gate>
<gate>
<ID>50</ID>
<type>DE_TO</type>
<position>236,35</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a6</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_AND2</type>
<position>231,86</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND2</type>
<position>231,82</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_OR4</type>
<position>237.5,89</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>29 </input>
<input>
<ID>IN_2</ID>22 </input>
<input>
<ID>IN_3</ID>21 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>54</ID>
<type>DE_TO</type>
<position>243.5,89</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a1</lparam></gate>
<gate>
<ID>56</ID>
<type>AE_FULLADDER_4BIT</type>
<position>78.5,-32</position>
<input>
<ID>IN_3</ID>199 </input>
<input>
<ID>IN_B_0</ID>199 </input>
<input>
<ID>IN_B_1</ID>110 </input>
<input>
<ID>IN_B_2</ID>106 </input>
<input>
<ID>IN_B_3</ID>85 </input>
<output>
<ID>OUT_0</ID>202 </output>
<output>
<ID>OUT_1</ID>200 </output>
<output>
<ID>OUT_2</ID>201 </output>
<output>
<ID>OUT_3</ID>203 </output>
<output>
<ID>carry_out</ID>60 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>57</ID>
<type>AE_FULLADDER_4BIT</type>
<position>78.5,-48</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>106 </input>
<input>
<ID>IN_2</ID>85 </input>
<output>
<ID>OUT_0</ID>229 </output>
<output>
<ID>OUT_1</ID>207 </output>
<output>
<ID>OUT_2</ID>206 </output>
<output>
<ID>OUT_3</ID>205 </output>
<input>
<ID>carry_in</ID>60 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_FULLADDER_4BIT</type>
<position>112,-13</position>
<input>
<ID>IN_2</ID>202 </input>
<input>
<ID>IN_3</ID>200 </input>
<input>
<ID>IN_B_1</ID>202 </input>
<input>
<ID>IN_B_2</ID>200 </input>
<input>
<ID>IN_B_3</ID>201 </input>
<output>
<ID>OUT_0</ID>214 </output>
<output>
<ID>OUT_1</ID>215 </output>
<output>
<ID>OUT_2</ID>216 </output>
<output>
<ID>OUT_3</ID>217 </output>
<output>
<ID>carry_out</ID>210 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_FULLADDER_4BIT</type>
<position>112,-29</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>203 </input>
<input>
<ID>IN_2</ID>229 </input>
<input>
<ID>IN_3</ID>207 </input>
<input>
<ID>IN_B_0</ID>203 </input>
<input>
<ID>IN_B_1</ID>229 </input>
<input>
<ID>IN_B_2</ID>207 </input>
<input>
<ID>IN_B_3</ID>206 </input>
<output>
<ID>OUT_0</ID>218 </output>
<output>
<ID>OUT_1</ID>219 </output>
<output>
<ID>OUT_2</ID>220 </output>
<output>
<ID>OUT_3</ID>221 </output>
<input>
<ID>carry_in</ID>210 </input>
<output>
<ID>carry_out</ID>212 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_FULLADDER_4BIT</type>
<position>112,-45</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>205 </input>
<input>
<ID>IN_B_0</ID>205 </input>
<output>
<ID>OUT_0</ID>222 </output>
<output>
<ID>OUT_1</ID>223 </output>
<output>
<ID>OUT_2</ID>224 </output>
<output>
<ID>OUT_3</ID>225 </output>
<input>
<ID>carry_in</ID>212 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,85</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>65</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>44,-23.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>41 </input>
<input>
<ID>IN_3</ID>40 </input>
<output>
<ID>OUT_0</ID>59 </output>
<output>
<ID>OUT_1</ID>55 </output>
<output>
<ID>OUT_2</ID>54 </output>
<output>
<ID>OUT_3</ID>53 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>66</ID>
<type>DE_OR8</type>
<position>31.5,-34.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>35 </input>
<input>
<ID>IN_3</ID>34 </input>
<input>
<ID>IN_4</ID>30 </input>
<input>
<ID>IN_5</ID>31 </input>
<input>
<ID>IN_6</ID>32 </input>
<input>
<ID>IN_7</ID>33 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>67</ID>
<type>FF_GND</type>
<position>27.5,-33</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_OR2</type>
<position>31.5,-12.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_OR4</type>
<position>31.5,-26.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>31 </input>
<input>
<ID>IN_3</ID>38 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>70</ID>
<type>AE_OR4</type>
<position>31.5,-18.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>32 </input>
<input>
<ID>IN_3</ID>43 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_OR4</type>
<position>45,-11.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>37 </input>
<input>
<ID>IN_3</ID>36 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_OR2</type>
<position>53,-3.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>BB_CLOCK</type>
<position>46,-46</position>
<output>
<ID>CLK</ID>61 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>52.5,-44</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_REGISTER4</type>
<position>52.5,-31.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>54 </input>
<input>
<ID>IN_3</ID>53 </input>
<output>
<ID>OUT_0</ID>199 </output>
<output>
<ID>OUT_1</ID>110 </output>
<output>
<ID>OUT_2</ID>106 </output>
<output>
<ID>OUT_3</ID>85 </output>
<input>
<ID>clear</ID>107 </input>
<input>
<ID>clock</ID>61 </input>
<input>
<ID>load</ID>58 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>79</ID>
<type>AE_SMALL_INVERTER</type>
<position>226,81</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>80</ID>
<type>BM_NORX2</type>
<position>231,90</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_AND2</type>
<position>227,61</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AE_OR4</type>
<position>238,53</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>44 </input>
<input>
<ID>IN_2</ID>46 </input>
<input>
<ID>IN_3</ID>47 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_AND2</type>
<position>231,56</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_AND2</type>
<position>231,52</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>HA_JUNC_2</type>
<position>166,49.5</position>
<input>
<ID>N_in0</ID>111 </input>
<input>
<ID>N_in1</ID>26 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>HA_JUNC_2</type>
<position>166,50.5</position>
<input>
<ID>N_in0</ID>112 </input>
<input>
<ID>N_in1</ID>28 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>HA_JUNC_2</type>
<position>166,51.5</position>
<input>
<ID>N_in0</ID>113 </input>
<input>
<ID>N_in1</ID>27 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>HA_JUNC_2</type>
<position>166,52.5</position>
<input>
<ID>N_in0</ID>114 </input>
<input>
<ID>N_in1</ID>23 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>CC_PULSE</type>
<position>-4,-7</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>90</ID>
<type>CC_PULSE</type>
<position>0,15.5</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>91</ID>
<type>CC_PULSE</type>
<position>-4,15.5</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>92</ID>
<type>CC_PULSE</type>
<position>-8,15.5</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>93</ID>
<type>CC_PULSE</type>
<position>0,8</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>94</ID>
<type>CC_PULSE</type>
<position>-4,8</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>95</ID>
<type>CC_PULSE</type>
<position>-8,8</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>96</ID>
<type>CC_PULSE</type>
<position>0,0.5</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>97</ID>
<type>CC_PULSE</type>
<position>-4,0.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>98</ID>
<type>CC_PULSE</type>
<position>-8,0.5</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>99</ID>
<type>DE_TO</type>
<position>-8,19.5</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t7</lparam></gate>
<gate>
<ID>100</ID>
<type>DE_TO</type>
<position>-4,19.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t8</lparam></gate>
<gate>
<ID>101</ID>
<type>DE_TO</type>
<position>0,19.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t9</lparam></gate>
<gate>
<ID>102</ID>
<type>DE_TO</type>
<position>-8,12</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t4</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>-4,12</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t5</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>0,12</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t6</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>-8,4.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t1</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>-4,4.5</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t2</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_TO</type>
<position>0,4.5</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t3</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>-4,-3</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID t0</lparam></gate>
<gate>
<ID>109</ID>
<type>CC_PULSE</type>
<position>-12,-10</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>-12,-6</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID tCE</lparam></gate>
<gate>
<ID>112</ID>
<type>AE_OR2</type>
<position>12,-6</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AE_OR2</type>
<position>12,-10</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_OR2</type>
<position>12,-14</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>102 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AE_OR2</type>
<position>12,-18</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>AE_OR2</type>
<position>12,-22</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_OR2</type>
<position>12,-26</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR2</type>
<position>12,-30</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>98 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_OR2</type>
<position>12,-34</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_OR2</type>
<position>12,-38</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_OR2</type>
<position>12,-42</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>7,-43</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t0</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>7,-37</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t1</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>7,-33</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t2</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>7,-29</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t3</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>7,-25</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t4</lparam></gate>
<gate>
<ID>129</ID>
<type>DA_FROM</type>
<position>7,-21</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t5</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>7,-17</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t6</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>7,-13</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t7</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>7,-9</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t8</lparam></gate>
<gate>
<ID>133</ID>
<type>DA_FROM</type>
<position>7,-5</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID t9</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>7,-41</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>7,-39</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>7,-35</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>137</ID>
<type>DA_FROM</type>
<position>7,-31</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>138</ID>
<type>DA_FROM</type>
<position>7,-27</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>139</ID>
<type>DA_FROM</type>
<position>7,-23</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>140</ID>
<type>DA_FROM</type>
<position>7,-19</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>141</ID>
<type>DA_FROM</type>
<position>7,-15</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>7,-11</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>7,-7</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>144</ID>
<type>DA_FROM</type>
<position>54.5,-44</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID tCE</lparam></gate>
<gate>
<ID>145</ID>
<type>AE_OR2</type>
<position>53.5,-39</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>GA_LED</type>
<position>156.5,-12.5</position>
<input>
<ID>N_in0</ID>214 </input>
<input>
<ID>N_in1</ID>111 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>156.5,-15.5</position>
<input>
<ID>N_in0</ID>215 </input>
<input>
<ID>N_in1</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>156.5,-18.5</position>
<input>
<ID>N_in0</ID>216 </input>
<input>
<ID>N_in1</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>GA_LED</type>
<position>156.5,-21.5</position>
<input>
<ID>N_in0</ID>217 </input>
<input>
<ID>N_in1</ID>114 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>GA_LED</type>
<position>156.5,-26.5</position>
<input>
<ID>N_in0</ID>218 </input>
<input>
<ID>N_in1</ID>191 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>GA_LED</type>
<position>156.5,-29.5</position>
<input>
<ID>N_in0</ID>219 </input>
<input>
<ID>N_in1</ID>192 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>GA_LED</type>
<position>156.5,-32.5</position>
<input>
<ID>N_in0</ID>220 </input>
<input>
<ID>N_in1</ID>193 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>156.5,-35.5</position>
<input>
<ID>N_in0</ID>221 </input>
<input>
<ID>N_in1</ID>194 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>GA_LED</type>
<position>156.5,-39.5</position>
<input>
<ID>N_in0</ID>222 </input>
<input>
<ID>N_in1</ID>195 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>156.5,-42.5</position>
<input>
<ID>N_in0</ID>223 </input>
<input>
<ID>N_in1</ID>196 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>GA_LED</type>
<position>156.5,-45.5</position>
<input>
<ID>N_in0</ID>224 </input>
<input>
<ID>N_in1</ID>197 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>156.5,-48.5</position>
<input>
<ID>N_in0</ID>225 </input>
<input>
<ID>N_in1</ID>198 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>BM_NORX2</type>
<position>233,-50</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>AE_OR3</type>
<position>235,-14</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>118 </input>
<input>
<ID>IN_2</ID>117 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>163</ID>
<type>AE_SMALL_INVERTER</type>
<position>230,-12</position>
<input>
<ID>IN_0</ID>131 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>164</ID>
<type>BM_NORX2</type>
<position>229,-15</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>AE_SMALL_INVERTER</type>
<position>228,-23</position>
<input>
<ID>IN_0</ID>131 </input>
<output>
<ID>OUT_0</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_AND3</type>
<position>233,-63</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>123 </input>
<input>
<ID>IN_2</ID>130 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>167</ID>
<type>AE_SMALL_INVERTER</type>
<position>228,-29</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>168</ID>
<type>AE_SMALL_INVERTER</type>
<position>228,-33</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>169</ID>
<type>AE_OR2</type>
<position>239,-37</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND2</type>
<position>233,-40</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>BM_NORX2</type>
<position>233,-36</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AE_SMALL_INVERTER</type>
<position>228,-41</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>173</ID>
<type>AE_OR3</type>
<position>233,-45</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>131 </input>
<input>
<ID>IN_2</ID>130 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>174</ID>
<type>AE_SMALL_INVERTER</type>
<position>228,-43</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>175</ID>
<type>AE_OR4</type>
<position>240,-55</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>120 </input>
<input>
<ID>IN_2</ID>121 </input>
<input>
<ID>IN_3</ID>122 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_AND2</type>
<position>233,-54</position>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_AND2</type>
<position>233,-58</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>149 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>AE_SMALL_INVERTER</type>
<position>228,-53</position>
<input>
<ID>IN_0</ID>131 </input>
<output>
<ID>OUT_0</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>179</ID>
<type>AE_SMALL_INVERTER</type>
<position>228,-59</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>180</ID>
<type>AE_OR4</type>
<position>234.5,-4</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>127 </input>
<input>
<ID>IN_2</ID>151 </input>
<input>
<ID>IN_3</ID>152 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>181</ID>
<type>BM_NORX2</type>
<position>228.5,-5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_AND2</type>
<position>228.5,-9</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>AE_SMALL_INVERTER</type>
<position>228,-63</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_AND2</type>
<position>233,-32</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>139 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>185</ID>
<type>DE_TO</type>
<position>240.5,-4</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b2</lparam></gate>
<gate>
<ID>186</ID>
<type>DE_TO</type>
<position>240,-14</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b3</lparam></gate>
<gate>
<ID>187</ID>
<type>DE_TO</type>
<position>246,-27</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b4</lparam></gate>
<gate>
<ID>188</ID>
<type>DE_TO</type>
<position>244,-37</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b5</lparam></gate>
<gate>
<ID>189</ID>
<type>DE_TO</type>
<position>246,-55</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b7</lparam></gate>
<gate>
<ID>190</ID>
<type>DE_TO</type>
<position>238,-45</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b6</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_AND2</type>
<position>233,6</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_AND2</type>
<position>233,2</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>193</ID>
<type>AE_OR4</type>
<position>239.5,9</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>133 </input>
<input>
<ID>IN_2</ID>126 </input>
<input>
<ID>IN_3</ID>125 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>194</ID>
<type>DE_TO</type>
<position>245.5,9</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b1</lparam></gate>
<gate>
<ID>195</ID>
<type>AE_SMALL_INVERTER</type>
<position>228,5</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>196</ID>
<type>AE_SMALL_INVERTER</type>
<position>228,1</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>197</ID>
<type>BM_NORX2</type>
<position>233,10</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND2</type>
<position>229,-19</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_OR4</type>
<position>240,-27</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>134 </input>
<input>
<ID>IN_2</ID>135 </input>
<input>
<ID>IN_3</ID>136 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_AND2</type>
<position>233,-24</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_AND2</type>
<position>233,-28</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>HA_JUNC_2</type>
<position>207,-26</position>
<input>
<ID>N_in0</ID>191 </input>
<input>
<ID>N_in1</ID>130 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>HA_JUNC_2</type>
<position>207,-25</position>
<input>
<ID>N_in0</ID>192 </input>
<input>
<ID>N_in1</ID>132 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>204</ID>
<type>HA_JUNC_2</type>
<position>207,-24</position>
<input>
<ID>N_in0</ID>193 </input>
<input>
<ID>N_in1</ID>131 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>HA_JUNC_2</type>
<position>207,-23</position>
<input>
<ID>N_in0</ID>194 </input>
<input>
<ID>N_in1</ID>127 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>BM_NORX2</type>
<position>233.5,-132.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>AE_OR3</type>
<position>235.5,-96.5</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>156 </input>
<input>
<ID>IN_2</ID>155 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>208</ID>
<type>AE_SMALL_INVERTER</type>
<position>230.5,-94.5</position>
<input>
<ID>IN_0</ID>169 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>209</ID>
<type>BM_NORX2</type>
<position>229.5,-97.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>AE_SMALL_INVERTER</type>
<position>228.5,-105.5</position>
<input>
<ID>IN_0</ID>169 </input>
<output>
<ID>OUT_0</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_AND3</type>
<position>233.5,-145.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>161 </input>
<input>
<ID>IN_2</ID>168 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>212</ID>
<type>AE_SMALL_INVERTER</type>
<position>228.5,-111.5</position>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>213</ID>
<type>AE_SMALL_INVERTER</type>
<position>228.5,-115.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>214</ID>
<type>AE_OR2</type>
<position>239.5,-119.5</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>180 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_AND2</type>
<position>233.5,-122.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>182 </input>
<output>
<ID>OUT</ID>180 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>BM_NORX2</type>
<position>233.5,-118.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>AE_SMALL_INVERTER</type>
<position>228.5,-123.5</position>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>182 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>218</ID>
<type>AE_OR3</type>
<position>233.5,-127.5</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>169 </input>
<input>
<ID>IN_2</ID>168 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>219</ID>
<type>AE_SMALL_INVERTER</type>
<position>228.5,-125.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>184 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>220</ID>
<type>AE_OR4</type>
<position>240.5,-137.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>158 </input>
<input>
<ID>IN_2</ID>159 </input>
<input>
<ID>IN_3</ID>160 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>233.5,-136.5</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_AND2</type>
<position>233.5,-140.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>223</ID>
<type>AE_SMALL_INVERTER</type>
<position>228.5,-135.5</position>
<input>
<ID>IN_0</ID>169 </input>
<output>
<ID>OUT_0</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>224</ID>
<type>AE_SMALL_INVERTER</type>
<position>228.5,-141.5</position>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>225</ID>
<type>AE_OR4</type>
<position>235,-86.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>165 </input>
<input>
<ID>IN_2</ID>189 </input>
<input>
<ID>IN_3</ID>190 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>226</ID>
<type>BM_NORX2</type>
<position>229,-87.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_AND2</type>
<position>229,-91.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AE_SMALL_INVERTER</type>
<position>228.5,-145.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_AND2</type>
<position>233.5,-114.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>177 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>DE_TO</type>
<position>241.5,-86.5</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c2</lparam></gate>
<gate>
<ID>231</ID>
<type>DE_TO</type>
<position>240.5,-96.5</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c3</lparam></gate>
<gate>
<ID>232</ID>
<type>DE_TO</type>
<position>246.5,-109.5</position>
<input>
<ID>IN_0</ID>178 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c4</lparam></gate>
<gate>
<ID>233</ID>
<type>DE_TO</type>
<position>244.5,-119.5</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c5</lparam></gate>
<gate>
<ID>234</ID>
<type>DE_TO</type>
<position>246.5,-137.5</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c7</lparam></gate>
<gate>
<ID>235</ID>
<type>DE_TO</type>
<position>238.5,-127.5</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c6</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>233.5,-76.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>166 </input>
<output>
<ID>OUT</ID>164 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>AA_AND2</type>
<position>233.5,-80.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>167 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>238</ID>
<type>AE_OR4</type>
<position>240,-73.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>171 </input>
<input>
<ID>IN_2</ID>164 </input>
<input>
<ID>IN_3</ID>163 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>239</ID>
<type>DE_TO</type>
<position>246,-73.5</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c1</lparam></gate>
<gate>
<ID>240</ID>
<type>AE_SMALL_INVERTER</type>
<position>228.5,-77.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_SMALL_INVERTER</type>
<position>228.5,-81.5</position>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>167 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>242</ID>
<type>BM_NORX2</type>
<position>233.5,-72.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_AND2</type>
<position>229.5,-101.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>AE_OR4</type>
<position>240.5,-109.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>172 </input>
<input>
<ID>IN_2</ID>173 </input>
<input>
<ID>IN_3</ID>174 </input>
<output>
<ID>OUT</ID>178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>245</ID>
<type>AA_AND2</type>
<position>233.5,-106.5</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_AND2</type>
<position>233.5,-110.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>176 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>247</ID>
<type>HA_JUNC_2</type>
<position>207.5,-108.5</position>
<input>
<ID>N_in0</ID>195 </input>
<input>
<ID>N_in1</ID>168 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>HA_JUNC_2</type>
<position>207.5,-107.5</position>
<input>
<ID>N_in0</ID>196 </input>
<input>
<ID>N_in1</ID>170 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>249</ID>
<type>HA_JUNC_2</type>
<position>207.5,-106.5</position>
<input>
<ID>N_in0</ID>197 </input>
<input>
<ID>N_in1</ID>169 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>HA_JUNC_2</type>
<position>207.5,-105.5</position>
<input>
<ID>N_in0</ID>198 </input>
<input>
<ID>N_in1</ID>165 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>97.5,-55</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>207 </input>
<input>
<ID>IN_2</ID>206 </input>
<input>
<ID>IN_3</ID>205 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>254</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>100.5,-4</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>200 </input>
<input>
<ID>IN_2</ID>201 </input>
<input>
<ID>IN_3</ID>203 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_LABEL</type>
<position>162,-12</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>259</ID>
<type>AA_LABEL</type>
<position>162,-15</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>AA_LABEL</type>
<position>162,-17.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>AA_LABEL</type>
<position>162,-20.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>160,-25.5</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>263</ID>
<type>AA_LABEL</type>
<position>159.5,-28.5</position>
<gparam>LABEL_TEXT 5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>159.5,-32</position>
<gparam>LABEL_TEXT 6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>265</ID>
<type>AA_LABEL</type>
<position>159.5,-35</position>
<gparam>LABEL_TEXT 7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>266</ID>
<type>AA_LABEL</type>
<position>160,-39</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>AA_LABEL</type>
<position>160,-42</position>
<gparam>LABEL_TEXT 9</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>268</ID>
<type>AA_LABEL</type>
<position>160,-44.5</position>
<gparam>LABEL_TEXT 10</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>AA_LABEL</type>
<position>160.5,-48</position>
<gparam>LABEL_TEXT 11</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>271</ID>
<type>AA_LABEL</type>
<position>162,-7.5</position>
<gparam>LABEL_TEXT 2 do potegi</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>273</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>177.5,-17</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>114 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 8</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>274</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>175,-31</position>
<input>
<ID>IN_0</ID>191 </input>
<input>
<ID>IN_1</ID>192 </input>
<input>
<ID>IN_2</ID>193 </input>
<input>
<ID>IN_3</ID>194 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 13</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,66,236,66</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,68,230,68</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,61,230,64</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,65,230,66</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,28,235,30</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,30,235,30</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234,26,235,26</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<connection>
<GID>16</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,22,234,24</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,24,235,24</points>
<connection>
<GID>15</GID>
<name>IN_2</name></connection>
<intersection>234 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,17,235,22</points>
<connection>
<GID>15</GID>
<name>IN_3</name></connection>
<intersection>17 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>234,17,235,17</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,17,228,17</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>241.5,89,241.5,89</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<connection>
<GID>54</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,82,234.5,86</points>
<connection>
<GID>53</GID>
<name>IN_3</name></connection>
<intersection>82 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>234,82,234.5,82</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,86,234,88</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,88,234.5,88</points>
<connection>
<GID>53</GID>
<name>IN_2</name></connection>
<intersection>234 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,52.5,173,92</points>
<intersection>52.5 2</intersection>
<intersection>77 6</intersection>
<intersection>92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173,92,234.5,92</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167,52.5,196,52.5</points>
<connection>
<GID>88</GID>
<name>N_in1</name></connection>
<intersection>173 0</intersection>
<intersection>196 21</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>173,77,229.5,77</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>173 0</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>196,52.5,196,56</points>
<intersection>52.5 2</intersection>
<intersection>56 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>196,56,235,56</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>196 21</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,85,228,85</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>228,81,228,81</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172.5,51,224,51</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>172.5 50</intersection>
<intersection>185 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>185,15,185,89</points>
<intersection>15 47</intersection>
<intersection>21 64</intersection>
<intersection>29 40</intersection>
<intersection>33 22</intersection>
<intersection>39 63</intersection>
<intersection>43 18</intersection>
<intersection>51 1</intersection>
<intersection>60 66</intersection>
<intersection>64 62</intersection>
<intersection>70 28</intersection>
<intersection>74 38</intersection>
<intersection>81 65</intersection>
<intersection>89 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>185,89,228,89</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>185 5</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>185,43,228,43</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>185 5</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>185,33,228,33</points>
<connection>
<GID>13</GID>
<name>IN_2</name></connection>
<intersection>185 5</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>185,70,223.5,70</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>185 5</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>185,74,223.5,74</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>185 5</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>185,29,228,29</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>185 5</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>185,15,228,15</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>185 5</intersection></hsegment>
<vsegment>
<ID>50</ID>
<points>172.5,49.5,172.5,51</points>
<intersection>49.5 51</intersection>
<intersection>51 1</intersection></vsegment>
<hsegment>
<ID>51</ID>
<points>167,49.5,172.5,49.5</points>
<connection>
<GID>85</GID>
<name>N_in1</name></connection>
<intersection>172.5 50</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>185,64,224,64</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>185 5</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>185,39,224,39</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>185 5</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>185,21,224,21</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>185 5</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>185,81,224,81</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>185 5</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>185,60,224,60</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>185 5</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,19,176,87</points>
<intersection>19 41</intersection>
<intersection>27 37</intersection>
<intersection>31 35</intersection>
<intersection>35 17</intersection>
<intersection>45 30</intersection>
<intersection>49 15</intersection>
<intersection>51.5 45</intersection>
<intersection>57 5</intersection>
<intersection>68 39</intersection>
<intersection>72 25</intersection>
<intersection>76 11</intersection>
<intersection>83 1</intersection>
<intersection>87 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,83,228,83</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>176,87,228,87</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>176,57,224,57</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>176,76,223.5,76</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>176,49,228,49</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>176,35,228,35</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>176,72,223.5,72</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>176,45,228,45</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>176,31,228,31</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>176,27,224,27</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>176,68,226,68</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>176,19,228,19</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>167,51.5,176,51.5</points>
<connection>
<GID>87</GID>
<name>N_in1</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181,17,181,91</points>
<intersection>17 33</intersection>
<intersection>23 28</intersection>
<intersection>25 18</intersection>
<intersection>37 16</intersection>
<intersection>41 25</intersection>
<intersection>47 12</intersection>
<intersection>55 8</intersection>
<intersection>62 26</intersection>
<intersection>66 31</intersection>
<intersection>79 1</intersection>
<intersection>85 2</intersection>
<intersection>91 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171.5,79,229.5,79</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>171.5 36</intersection>
<intersection>181 0</intersection>
<intersection>189 38</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>181,85,224,85</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>181,91,228,91</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>167,55,228,55</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>167 45</intersection>
<intersection>171.5 36</intersection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>181,47,224,47</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>181,37,224,37</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>181,25,228,25</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>181,41,228,41</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>181,62,224,62</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>181,23,228,23</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>181,66,224,66</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>181,17,224,17</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>171.5,55,171.5,79</points>
<intersection>55 8</intersection>
<intersection>79 1</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>189,53,189,79</points>
<intersection>53 46</intersection>
<intersection>79 1</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>167,50.5,167,55</points>
<connection>
<GID>86</GID>
<name>N_in1</name></connection>
<intersection>55 8</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>189,53,228,53</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>189 38</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234,90,234.5,90</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<connection>
<GID>80</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>15,-38,28.5,-38</points>
<connection>
<GID>66</GID>
<name>IN_4</name></connection>
<connection>
<GID>120</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-37,24,-27.5</points>
<intersection>-37 2</intersection>
<intersection>-30 4</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24,-37,28.5,-37</points>
<connection>
<GID>66</GID>
<name>IN_5</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24,-27.5,28.5,-27.5</points>
<connection>
<GID>69</GID>
<name>IN_2</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>15,-30,24,-30</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-36,24.5,-19.5</points>
<intersection>-36 2</intersection>
<intersection>-22.5 1</intersection>
<intersection>-19.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-22.5,24.5,-22.5</points>
<intersection>15 4</intersection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-36,28.5,-36</points>
<connection>
<GID>66</GID>
<name>IN_6</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24.5,-19.5,28.5,-19.5</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>24.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-22.5,15,-22</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>-22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-35,25,-15.5</points>
<intersection>-35 2</intersection>
<intersection>-23.5 3</intersection>
<intersection>-18.5 1</intersection>
<intersection>-15.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-18.5,25,-18.5</points>
<intersection>15 5</intersection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-35,28.5,-35</points>
<connection>
<GID>66</GID>
<name>IN_7</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25,-23.5,28.5,-23.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>25,-15.5,28.5,-15.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>15,-18.5,15,-14</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-34,25.5,-6</points>
<intersection>-34 2</intersection>
<intersection>-11.5 3</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-6,25.5,-6</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-34,28.5,-34</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25.5,-11.5,28.5,-11.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-33,28.5,-31</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-34.5,37,-14.5</points>
<intersection>-34.5 8</intersection>
<intersection>-24.5 4</intersection>
<intersection>-14.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37,-24.5,41,-24.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>37,-14.5,42,-14.5</points>
<connection>
<GID>72</GID>
<name>IN_3</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>35.5,-34.5,37,-34.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-26.5,36.5,-12.5</points>
<intersection>-26.5 2</intersection>
<intersection>-23.5 1</intersection>
<intersection>-12.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-23.5,41,-23.5</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-26.5,36.5,-26.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36.5,-12.5,42,-12.5</points>
<connection>
<GID>72</GID>
<name>IN_2</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-29.5,24,-28.5</points>
<intersection>-29.5 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-28.5,24,-28.5</points>
<intersection>20.5 3</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-29.5,28.5,-29.5</points>
<connection>
<GID>69</GID>
<name>IN_3</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20.5,-34,20.5,-28.5</points>
<intersection>-34 4</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>15,-34,20.5,-34</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>20.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-25.5,24,-17.5</points>
<intersection>-25.5 2</intersection>
<intersection>-20.5 1</intersection>
<intersection>-17.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-20.5,24,-20.5</points>
<intersection>15 4</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-25.5,28.5,-25.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24,-17.5,28.5,-17.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-20.5,15,-18</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-21.5,38,-12.5</points>
<intersection>-21.5 3</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-12.5,38,-12.5</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38,-21.5,41,-21.5</points>
<connection>
<GID>65</GID>
<name>IN_3</name></connection>
<intersection>38 0</intersection>
<intersection>40 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>40,-21.5,40,-8.5</points>
<intersection>-21.5 3</intersection>
<intersection>-8.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>40,-8.5,42,-8.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>40 6</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-22.5,36.5,-18.5</points>
<intersection>-22.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-22.5,41,-22.5</points>
<connection>
<GID>65</GID>
<name>IN_2</name></connection>
<intersection>36.5 0</intersection>
<intersection>39 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-18.5,36.5,-18.5</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>39,-22.5,39,-10.5</points>
<intersection>-22.5 1</intersection>
<intersection>-10.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>39,-10.5,42,-10.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>39 5</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-16.5,24.5,-13.5</points>
<intersection>-16.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-16.5,24.5,-16.5</points>
<intersection>15 3</intersection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-13.5,28.5,-13.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,-16.5,15,-10</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>-16.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-24.5,24,-21.5</points>
<intersection>-24.5 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-24.5,24,-24.5</points>
<intersection>15 3</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-21.5,28.5,-21.5</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,-26,15,-24.5</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,54,234,56</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>234,54,235,54</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>234 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-42,22,-4.5</points>
<intersection>-42 4</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22,-4.5,50,-4.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>15,-42,22,-42</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234,52,235,52</points>
<connection>
<GID>82</GID>
<name>IN_2</name></connection>
<connection>
<GID>84</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,48,234.5,50</points>
<intersection>48 1</intersection>
<intersection>50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,48,234.5,48</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234.5,50,235,50</points>
<connection>
<GID>82</GID>
<name>IN_3</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,57,228,57</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<connection>
<GID>83</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,51,228,51</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,47,228,47</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,53,242,53</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>82</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,43,240,43</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-29.5,42.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_3</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-29.5,48.5,-29.5</points>
<connection>
<GID>76</GID>
<name>IN_3</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-30.5,43.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_2</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-30.5,48.5,-30.5</points>
<connection>
<GID>76</GID>
<name>IN_2</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-31.5,44.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_1</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-31.5,48.5,-31.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,40,234,42</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<connection>
<GID>9</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-11.5,49,-2.5</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-2.5,50,-2.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-26.5,51.5,-15.5</points>
<connection>
<GID>76</GID>
<name>load</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-15.5,56,-15.5</points>
<intersection>51.5 0</intersection>
<intersection>56 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>56,-15.5,56,-3.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>-15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-32.5,45.5,-27.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-32.5,48.5,-32.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-40,77.5,-40</points>
<connection>
<GID>56</GID>
<name>carry_out</name></connection>
<connection>
<GID>57</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-42,46,-35.5</points>
<connection>
<GID>74</GID>
<name>CLK</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-35.5,51.5,-35.5</points>
<connection>
<GID>76</GID>
<name>clock</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,44,234,44</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>11</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,39,228,39</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,35,234,35</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<connection>
<GID>50</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,37,228,37</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,25,242,25</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<connection>
<GID>49</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,27,228,27</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,21,228,21</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,76,236.5,76</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,75,229.5,75</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<connection>
<GID>21</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,71,229.5,73</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-8,17.5,-8,17.5</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,17.5,-4,17.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.43359e-008,17.5,2.43359e-008,17.5</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,10,-8,10</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,10,-4,10</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<connection>
<GID>103</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-2.43359e-008,10,2.43359e-008,10</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<connection>
<GID>104</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,2.5,-8,2.5</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,2.5,-4,2.5</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.43359e-008,2.5,2.43359e-008,2.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<connection>
<GID>107</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-5,-4,-5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-8,-12,-8</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-43,9,-43</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<connection>
<GID>123</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-25,72.5,-25</points>
<intersection>56.5 11</intersection>
<intersection>72.5 12</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>56.5,-29.5,56.5,-25</points>
<connection>
<GID>76</GID>
<name>OUT_3</name></connection>
<intersection>-25 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>72.5,-30,72.5,-25</points>
<intersection>-30 13</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>61,-30,74.5,-30</points>
<connection>
<GID>56</GID>
<name>IN_B_3</name></connection>
<intersection>61 14</intersection>
<intersection>72.5 12</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>61,-52,61,-30</points>
<intersection>-52 15</intersection>
<intersection>-30 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>61,-52,74.5,-52</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<intersection>61 14</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-37,9,-37</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<connection>
<GID>125</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-33,9,-33</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<connection>
<GID>126</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-29,9,-29</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-25,9,-25</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<connection>
<GID>128</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-21,9,-21</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-17,9,-17</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-13,9,-13</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<connection>
<GID>131</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-9,9,-9</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<connection>
<GID>132</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-5,9,-5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-41,9,-41</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-39,9,-39</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<connection>
<GID>135</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-35,9,-35</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<connection>
<GID>136</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-31,9,-31</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<connection>
<GID>137</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-27,9,-27</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-23,9,-23</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-19,9,-19</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-15,9,-15</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-11,9,-11</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<connection>
<GID>142</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-7,9,-7</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<connection>
<GID>143</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-30.5,57.5,-29</points>
<intersection>-30.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-29,74.5,-29</points>
<connection>
<GID>56</GID>
<name>IN_B_2</name></connection>
<intersection>57.5 0</intersection>
<intersection>68.5 13</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-30.5,57.5,-30.5</points>
<connection>
<GID>76</GID>
<name>OUT_2</name></connection>
<intersection>57.5 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>68.5,-51,68.5,-29</points>
<intersection>-51 14</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>68.5,-51,74.5,-51</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>68.5 13</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>53.5,-36,53.5,-35.5</points>
<connection>
<GID>76</GID>
<name>clear</name></connection>
<connection>
<GID>145</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>54.5,-42,54.5,-42</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<connection>
<GID>145</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>52.5,-42,52.5,-42</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<connection>
<GID>145</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-50,63,-28</points>
<intersection>-50 9</intersection>
<intersection>-31.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-31.5,63,-31.5</points>
<connection>
<GID>76</GID>
<name>OUT_1</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-28,74.5,-28</points>
<connection>
<GID>56</GID>
<name>IN_B_1</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>63,-50,74.5,-50</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-18,158,49.5</points>
<intersection>-18 3</intersection>
<intersection>-12.5 2</intersection>
<intersection>49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158,49.5,165,49.5</points>
<connection>
<GID>85</GID>
<name>N_in0</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-12.5,158,-12.5</points>
<connection>
<GID>147</GID>
<name>N_in1</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>158,-18,174.5,-18</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,-17,158.5,50.5</points>
<intersection>-17 3</intersection>
<intersection>-15.5 2</intersection>
<intersection>50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158.5,50.5,165,50.5</points>
<connection>
<GID>86</GID>
<name>N_in0</name></connection>
<intersection>158.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-15.5,158.5,-15.5</points>
<connection>
<GID>148</GID>
<name>N_in1</name></connection>
<intersection>158.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>158.5,-17,174.5,-17</points>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<intersection>158.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159.5,-18.5,159.5,51.5</points>
<intersection>-18.5 2</intersection>
<intersection>-16 3</intersection>
<intersection>51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>159.5,51.5,165,51.5</points>
<connection>
<GID>87</GID>
<name>N_in0</name></connection>
<intersection>159.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-18.5,159.5,-18.5</points>
<connection>
<GID>149</GID>
<name>N_in1</name></connection>
<intersection>159.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>159.5,-16,174.5,-16</points>
<connection>
<GID>273</GID>
<name>IN_2</name></connection>
<intersection>159.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160.5,-21.5,160.5,52.5</points>
<intersection>-21.5 2</intersection>
<intersection>-15 3</intersection>
<intersection>52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160.5,52.5,165,52.5</points>
<connection>
<GID>88</GID>
<name>N_in0</name></connection>
<intersection>160.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-21.5,160.5,-21.5</points>
<connection>
<GID>150</GID>
<name>N_in1</name></connection>
<intersection>160.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>160.5,-15,174.5,-15</points>
<connection>
<GID>273</GID>
<name>IN_3</name></connection>
<intersection>160.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-14,238,-14</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232,-12,232,-12</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232,-19,232,-16</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<connection>
<GID>162</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232,-15,232,-14</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<connection>
<GID>162</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,-52,237,-50</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236,-50,237,-50</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>237 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,-54,237,-54</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<connection>
<GID>176</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-58,236,-56</points>
<connection>
<GID>177</GID>
<name>OUT</name></connection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236,-56,237,-56</points>
<connection>
<GID>175</GID>
<name>IN_2</name></connection>
<intersection>236 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,-63,237,-58</points>
<connection>
<GID>175</GID>
<name>IN_3</name></connection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>236,-63,237,-63</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<intersection>237 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-63,230,-63</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>243.5,9,243.5,9</points>
<connection>
<GID>193</GID>
<name>OUT</name></connection>
<connection>
<GID>194</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,2,236.5,6</points>
<connection>
<GID>193</GID>
<name>IN_3</name></connection>
<intersection>2 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>236,2,236.5,2</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<intersection>236.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,6,236,8</points>
<connection>
<GID>191</GID>
<name>OUT</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236,8,236.5,8</points>
<connection>
<GID>193</GID>
<name>IN_2</name></connection>
<intersection>236 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214,-23,214,12</points>
<intersection>-23 2</intersection>
<intersection>-3 6</intersection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214,12,236.5,12</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>208,-23,237,-23</points>
<connection>
<GID>205</GID>
<name>N_in1</name></connection>
<intersection>214 0</intersection>
<intersection>237 21</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>214,-3,231.5,-3</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>214 0</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>237,-24,237,-23</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>-23 2</intersection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,5,230,5</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>230,1,230,1</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213.5,-29,226,-29</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>213.5 50</intersection>
<intersection>226 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>226,-65,226,9</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>-65 47</intersection>
<intersection>-51 40</intersection>
<intersection>-47 22</intersection>
<intersection>-37 18</intersection>
<intersection>-29 1</intersection>
<intersection>-10 28</intersection>
<intersection>-6 38</intersection>
<intersection>9 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>226,9,230,9</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>226 5</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>226,-37,230,-37</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>226 5</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>226,-47,230,-47</points>
<connection>
<GID>173</GID>
<name>IN_2</name></connection>
<intersection>226 5</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>225.5,-10,226,-10</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>226 5</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>225.5,-6,226,-6</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>226 5</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>226,-51,230,-51</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>226 5</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>226,-65,230,-65</points>
<connection>
<GID>166</GID>
<name>IN_2</name></connection>
<intersection>226 5</intersection></hsegment>
<vsegment>
<ID>50</ID>
<points>213.5,-29,213.5,-26</points>
<intersection>-29 1</intersection>
<intersection>-26 51</intersection></vsegment>
<hsegment>
<ID>51</ID>
<points>208,-26,213.5,-26</points>
<connection>
<GID>202</GID>
<name>N_in1</name></connection>
<intersection>213.5 50</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217,-61,217,7</points>
<intersection>-61 41</intersection>
<intersection>-53 37</intersection>
<intersection>-49 35</intersection>
<intersection>-45 17</intersection>
<intersection>-35 30</intersection>
<intersection>-31 15</intersection>
<intersection>-24 45</intersection>
<intersection>-23 5</intersection>
<intersection>-12 39</intersection>
<intersection>-8 25</intersection>
<intersection>-4 11</intersection>
<intersection>3 1</intersection>
<intersection>7 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>217,3,230,3</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>217,7,230,7</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217,-23,226,-23</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>217,-4,225.5,-4</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>217,-31,230,-31</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>217,-45,230,-45</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>217,-8,225.5,-8</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>217,-35,230,-35</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>217,-49,230,-49</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>217,-53,226,-53</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>217,-12,228,-12</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>217,-61,230,-61</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>208,-24,217,-24</points>
<connection>
<GID>204</GID>
<name>N_in1</name></connection>
<intersection>217 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-63,222,11</points>
<intersection>-63 33</intersection>
<intersection>-57 28</intersection>
<intersection>-55 18</intersection>
<intersection>-43 16</intersection>
<intersection>-39 25</intersection>
<intersection>-33 12</intersection>
<intersection>-25 8</intersection>
<intersection>-18 26</intersection>
<intersection>-14 31</intersection>
<intersection>-1 1</intersection>
<intersection>5 2</intersection>
<intersection>11 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>212.5,-1,231.5,-1</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>212.5 36</intersection>
<intersection>222 0</intersection>
<intersection>230 38</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>222,5,226,5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>222,11,230,11</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>208,-25,230,-25</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<connection>
<GID>203</GID>
<name>N_in1</name></connection>
<intersection>212.5 36</intersection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>222,-33,226,-33</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>222,-43,226,-43</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>222,-55,230,-55</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>222,-39,230,-39</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>222,-18,226,-18</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>222,-57,230,-57</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>222,-14,226,-14</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>222,-63,226,-63</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>212.5,-25,212.5,-1</points>
<intersection>-25 8</intersection>
<intersection>-1 1</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>230,-27,230,-1</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,10,236.5,10</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<connection>
<GID>197</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-26,236,-24</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>236,-26,237,-26</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>236 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,-28,237,-28</points>
<connection>
<GID>199</GID>
<name>IN_2</name></connection>
<connection>
<GID>201</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,-32,236.5,-30</points>
<intersection>-32 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236,-32,236.5,-32</points>
<connection>
<GID>184</GID>
<name>OUT</name></connection>
<intersection>236.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>236.5,-30,237,-30</points>
<connection>
<GID>199</GID>
<name>IN_3</name></connection>
<intersection>236.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-23,230,-23</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<connection>
<GID>200</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-29,230,-29</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<connection>
<GID>201</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-33,230,-33</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<connection>
<GID>184</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-27,244,-27</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<connection>
<GID>199</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-37,242,-37</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<connection>
<GID>188</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-40,236,-38</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<connection>
<GID>169</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-36,236,-36</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<connection>
<GID>171</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-41,230,-41</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-45,236,-45</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<connection>
<GID>190</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-43,230,-43</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-55,244,-55</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<connection>
<GID>189</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-53,230,-53</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-59,230,-59</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-4,238.5,-4</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<connection>
<GID>185</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-5,231.5,-5</points>
<connection>
<GID>180</GID>
<name>IN_2</name></connection>
<connection>
<GID>181</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-9,231.5,-7</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<connection>
<GID>180</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-96.5,238.5,-96.5</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<connection>
<GID>231</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-94.5,232.5,-94.5</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-101.5,232.5,-98.5</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<connection>
<GID>207</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-97.5,232.5,-96.5</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<connection>
<GID>207</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-134.5,237.5,-132.5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>-132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236.5,-132.5,237.5,-132.5</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<intersection>237.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-136.5,237.5,-136.5</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<connection>
<GID>221</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,-140.5,236.5,-138.5</points>
<connection>
<GID>222</GID>
<name>OUT</name></connection>
<intersection>-138.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236.5,-138.5,237.5,-138.5</points>
<connection>
<GID>220</GID>
<name>IN_2</name></connection>
<intersection>236.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-145.5,237.5,-140.5</points>
<connection>
<GID>220</GID>
<name>IN_3</name></connection>
<intersection>-145.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>236.5,-145.5,237.5,-145.5</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>237.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-145.5,230.5,-145.5</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>244,-73.5,244,-73.5</points>
<connection>
<GID>238</GID>
<name>OUT</name></connection>
<connection>
<GID>239</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,-80.5,237,-76.5</points>
<connection>
<GID>238</GID>
<name>IN_3</name></connection>
<intersection>-80.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>236.5,-80.5,237,-80.5</points>
<connection>
<GID>237</GID>
<name>OUT</name></connection>
<intersection>237 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,-76.5,236.5,-74.5</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236.5,-74.5,237,-74.5</points>
<connection>
<GID>238</GID>
<name>IN_2</name></connection>
<intersection>236.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-105.5,214.5,-70.5</points>
<intersection>-105.5 2</intersection>
<intersection>-85.5 6</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214.5,-70.5,237,-70.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>214.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>208.5,-105.5,237.5,-105.5</points>
<connection>
<GID>250</GID>
<name>N_in1</name></connection>
<intersection>214.5 0</intersection>
<intersection>237.5 21</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>214.5,-85.5,232,-85.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>214.5 0</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>237.5,-106.5,237.5,-105.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>-105.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-77.5,230.5,-77.5</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>230.5,-81.5,230.5,-81.5</points>
<connection>
<GID>237</GID>
<name>IN_1</name></connection>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>214,-111.5,226.5,-111.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>214 50</intersection>
<intersection>226.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>226.5,-147.5,226.5,-73.5</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>-147.5 47</intersection>
<intersection>-133.5 40</intersection>
<intersection>-129.5 22</intersection>
<intersection>-119.5 18</intersection>
<intersection>-111.5 1</intersection>
<intersection>-92.5 28</intersection>
<intersection>-88.5 38</intersection>
<intersection>-73.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>226.5,-73.5,230.5,-73.5</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>226.5 5</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>226.5,-119.5,230.5,-119.5</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>226.5 5</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>226.5,-129.5,230.5,-129.5</points>
<connection>
<GID>218</GID>
<name>IN_2</name></connection>
<intersection>226.5 5</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>226,-92.5,226.5,-92.5</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<intersection>226.5 5</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>226,-88.5,226.5,-88.5</points>
<connection>
<GID>226</GID>
<name>IN_1</name></connection>
<intersection>226.5 5</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>226.5,-133.5,230.5,-133.5</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>226.5 5</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>226.5,-147.5,230.5,-147.5</points>
<connection>
<GID>211</GID>
<name>IN_2</name></connection>
<intersection>226.5 5</intersection></hsegment>
<vsegment>
<ID>50</ID>
<points>214,-111.5,214,-108.5</points>
<intersection>-111.5 1</intersection>
<intersection>-108.5 51</intersection></vsegment>
<hsegment>
<ID>51</ID>
<points>208.5,-108.5,214,-108.5</points>
<connection>
<GID>247</GID>
<name>N_in1</name></connection>
<intersection>214 50</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,-143.5,217.5,-75.5</points>
<intersection>-143.5 41</intersection>
<intersection>-135.5 37</intersection>
<intersection>-131.5 35</intersection>
<intersection>-127.5 17</intersection>
<intersection>-117.5 30</intersection>
<intersection>-113.5 15</intersection>
<intersection>-106.5 45</intersection>
<intersection>-105.5 5</intersection>
<intersection>-94.5 39</intersection>
<intersection>-90.5 25</intersection>
<intersection>-86.5 11</intersection>
<intersection>-79.5 1</intersection>
<intersection>-75.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>217.5,-79.5,230.5,-79.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>217.5,-75.5,230.5,-75.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217.5,-105.5,226.5,-105.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>217.5,-86.5,226,-86.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>217.5,-113.5,230.5,-113.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>217.5,-127.5,230.5,-127.5</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>217.5,-90.5,226,-90.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>217.5,-117.5,230.5,-117.5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>217.5,-131.5,230.5,-131.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>217.5,-135.5,226.5,-135.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>217.5,-94.5,228.5,-94.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>217.5,-143.5,230.5,-143.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>208.5,-106.5,217.5,-106.5</points>
<connection>
<GID>249</GID>
<name>N_in1</name></connection>
<intersection>217.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,-145.5,222.5,-71.5</points>
<intersection>-145.5 33</intersection>
<intersection>-139.5 28</intersection>
<intersection>-137.5 18</intersection>
<intersection>-125.5 16</intersection>
<intersection>-121.5 25</intersection>
<intersection>-115.5 12</intersection>
<intersection>-107.5 8</intersection>
<intersection>-100.5 26</intersection>
<intersection>-96.5 31</intersection>
<intersection>-83.5 1</intersection>
<intersection>-77.5 2</intersection>
<intersection>-71.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213,-83.5,232,-83.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>213 36</intersection>
<intersection>222.5 0</intersection>
<intersection>230.5 38</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>222.5,-77.5,226.5,-77.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>222.5,-71.5,230.5,-71.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>208.5,-107.5,230.5,-107.5</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<connection>
<GID>248</GID>
<name>N_in1</name></connection>
<intersection>213 36</intersection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>222.5,-115.5,226.5,-115.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>222.5,-125.5,226.5,-125.5</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>222.5,-137.5,230.5,-137.5</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>222.5,-121.5,230.5,-121.5</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>222.5,-100.5,226.5,-100.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>222.5,-139.5,230.5,-139.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>222.5,-96.5,226.5,-96.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>222.5,-145.5,226.5,-145.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>213,-107.5,213,-83.5</points>
<intersection>-107.5 8</intersection>
<intersection>-83.5 1</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>230.5,-109.5,230.5,-83.5</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>-83.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-72.5,237,-72.5</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<connection>
<GID>242</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,-108.5,236.5,-106.5</points>
<connection>
<GID>245</GID>
<name>OUT</name></connection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>236.5,-108.5,237.5,-108.5</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>236.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-110.5,237.5,-110.5</points>
<connection>
<GID>244</GID>
<name>IN_2</name></connection>
<connection>
<GID>246</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,-114.5,237,-112.5</points>
<intersection>-114.5 1</intersection>
<intersection>-112.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236.5,-114.5,237,-114.5</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<intersection>237 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237,-112.5,237.5,-112.5</points>
<connection>
<GID>244</GID>
<name>IN_3</name></connection>
<intersection>237 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-105.5,230.5,-105.5</points>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection>
<connection>
<GID>245</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-111.5,230.5,-111.5</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<connection>
<GID>246</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-115.5,230.5,-115.5</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<connection>
<GID>229</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244.5,-109.5,244.5,-109.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<connection>
<GID>244</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242.5,-119.5,242.5,-119.5</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<connection>
<GID>233</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,-122.5,236.5,-120.5</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<connection>
<GID>214</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,-118.5,236.5,-118.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<connection>
<GID>216</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-123.5,230.5,-123.5</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,-127.5,236.5,-127.5</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<connection>
<GID>235</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-125.5,230.5,-125.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>244.5,-137.5,244.5,-137.5</points>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<connection>
<GID>234</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-135.5,230.5,-135.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-141.5,230.5,-141.5</points>
<connection>
<GID>222</GID>
<name>IN_1</name></connection>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>239,-86.5,239.5,-86.5</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<connection>
<GID>230</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232,-87.5,232,-87.5</points>
<connection>
<GID>225</GID>
<name>IN_2</name></connection>
<connection>
<GID>226</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232,-91.5,232,-89.5</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<connection>
<GID>225</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-26.5,162,-26</points>
<intersection>-26.5 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-26.5,162,-26.5</points>
<connection>
<GID>151</GID>
<name>N_in1</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162,-26,206,-26</points>
<connection>
<GID>202</GID>
<name>N_in0</name></connection>
<intersection>162 0</intersection>
<intersection>164 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>164,-32,164,-26</points>
<intersection>-32 4</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>164,-32,172,-32</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>164 3</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157.5,-30.5,167,-30.5</points>
<intersection>157.5 3</intersection>
<intersection>164 4</intersection>
<intersection>167 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>167,-30.5,167,-25</points>
<intersection>-30.5 1</intersection>
<intersection>-25 6</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>157.5,-30.5,157.5,-29.5</points>
<connection>
<GID>152</GID>
<name>N_in1</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>164,-31,164,-30.5</points>
<intersection>-31 5</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>164,-31,172,-31</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>164 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>167,-25,206,-25</points>
<connection>
<GID>203</GID>
<name>N_in0</name></connection>
<intersection>167 2</intersection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-32.5,162,-24</points>
<intersection>-32.5 1</intersection>
<intersection>-30 3</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-32.5,162,-32.5</points>
<connection>
<GID>153</GID>
<name>N_in1</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162,-24,206,-24</points>
<connection>
<GID>204</GID>
<name>N_in0</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>162,-30,172,-30</points>
<connection>
<GID>274</GID>
<name>IN_2</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-35.5,163,-23</points>
<intersection>-35.5 1</intersection>
<intersection>-29 4</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-35.5,163,-35.5</points>
<connection>
<GID>154</GID>
<name>N_in1</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-23,206,-23</points>
<connection>
<GID>205</GID>
<name>N_in0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>163,-29,172,-29</points>
<connection>
<GID>274</GID>
<name>IN_3</name></connection>
<intersection>163 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-108.5,162.5,-39.5</points>
<intersection>-108.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-39.5,162.5,-39.5</points>
<connection>
<GID>155</GID>
<name>N_in1</name></connection>
<intersection>162.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-108.5,206.5,-108.5</points>
<connection>
<GID>247</GID>
<name>N_in0</name></connection>
<intersection>162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-107.5,162.5,-42.5</points>
<intersection>-107.5 1</intersection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-107.5,206.5,-107.5</points>
<connection>
<GID>248</GID>
<name>N_in0</name></connection>
<intersection>162.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-42.5,162.5,-42.5</points>
<connection>
<GID>156</GID>
<name>N_in1</name></connection>
<intersection>162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-106.5,162.5,-45.5</points>
<intersection>-106.5 2</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-45.5,162.5,-45.5</points>
<connection>
<GID>157</GID>
<name>N_in1</name></connection>
<intersection>162.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-106.5,206.5,-106.5</points>
<connection>
<GID>249</GID>
<name>N_in0</name></connection>
<intersection>162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-105.5,162.5,-48.5</points>
<intersection>-105.5 1</intersection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-105.5,206.5,-105.5</points>
<connection>
<GID>250</GID>
<name>N_in0</name></connection>
<intersection>162.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-48.5,162.5,-48.5</points>
<connection>
<GID>158</GID>
<name>N_in1</name></connection>
<intersection>162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-32.5,64,-27</points>
<intersection>-32.5 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-27,74.5,-27</points>
<connection>
<GID>56</GID>
<name>IN_B_0</name></connection>
<intersection>64 0</intersection>
<intersection>69 9</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-32.5,64,-32.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>69,-37,69,-27</points>
<intersection>-37 10</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>69,-37,74.5,-37</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>69 9</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-31.5,87.5,-31.5</points>
<connection>
<GID>56</GID>
<name>OUT_1</name></connection>
<intersection>87.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>87.5,-31.5,87.5,-4</points>
<intersection>-31.5 1</intersection>
<intersection>-10 6</intersection>
<intersection>-4 10</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>87.5,-10,108,-10</points>
<connection>
<GID>60</GID>
<name>IN_B_2</name></connection>
<intersection>87.5 5</intersection>
<intersection>102.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>102.5,-18,102.5,-10</points>
<intersection>-18 8</intersection>
<intersection>-10 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>102.5,-18,108,-18</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<intersection>102.5 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>87.5,-4,97.5,-4</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>87.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89,-31,108,-31</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>89 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89,-32.5,89,-3</points>
<intersection>-32.5 9</intersection>
<intersection>-31 1</intersection>
<intersection>-11 4</intersection>
<intersection>-3 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>89,-11,108,-11</points>
<connection>
<GID>60</GID>
<name>IN_B_3</name></connection>
<intersection>89 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>82.5,-32.5,89,-32.5</points>
<connection>
<GID>56</GID>
<name>OUT_2</name></connection>
<intersection>89 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>89,-3,97.5,-3</points>
<connection>
<GID>254</GID>
<name>IN_2</name></connection>
<intersection>89 3</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-30.5,86,-30.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>86 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>86,-30.5,86,-5</points>
<intersection>-30.5 1</intersection>
<intersection>-9 6</intersection>
<intersection>-5 10</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>86,-9,108,-9</points>
<connection>
<GID>60</GID>
<name>IN_B_1</name></connection>
<intersection>86 5</intersection>
<intersection>99.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>99.5,-17,99.5,-9</points>
<intersection>-17 8</intersection>
<intersection>-9 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>99.5,-17,108,-17</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>99.5 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>86,-5,97.5,-5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>86 5</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-33.5,89.5,-33.5</points>
<connection>
<GID>56</GID>
<name>OUT_3</name></connection>
<intersection>89.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>89.5,-33.5,89.5,-2</points>
<intersection>-33.5 1</intersection>
<intersection>-32 7</intersection>
<intersection>-24 5</intersection>
<intersection>-2 9</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>89.5,-24,108,-24</points>
<connection>
<GID>61</GID>
<name>IN_B_0</name></connection>
<intersection>89.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89.5,-32,108,-32</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>89.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>89.5,-2,97.5,-2</points>
<connection>
<GID>254</GID>
<name>IN_3</name></connection>
<intersection>89.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-49.5,101,-49.5</points>
<connection>
<GID>57</GID>
<name>OUT_3</name></connection>
<intersection>94.5 12</intersection>
<intersection>101 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>101,-49.5,101,-40</points>
<intersection>-49.5 1</intersection>
<intersection>-48 11</intersection>
<intersection>-40 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>101,-40,108,-40</points>
<connection>
<GID>62</GID>
<name>IN_B_0</name></connection>
<intersection>101 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>101,-48,108,-48</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>101 8</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>94.5,-53,94.5,-49.5</points>
<connection>
<GID>251</GID>
<name>IN_3</name></connection>
<intersection>-49.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-48.5,100.5,-48.5</points>
<connection>
<GID>57</GID>
<name>OUT_2</name></connection>
<intersection>92.5 12</intersection>
<intersection>100.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>100.5,-48.5,100.5,-27</points>
<intersection>-48.5 1</intersection>
<intersection>-47 11</intersection>
<intersection>-27 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>100.5,-27,108,-27</points>
<connection>
<GID>61</GID>
<name>IN_B_3</name></connection>
<intersection>100.5 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>100.5,-47,108,-47</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>100.5 8</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>92.5,-54,92.5,-48.5</points>
<intersection>-54 13</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>92.5,-54,94.5,-54</points>
<connection>
<GID>251</GID>
<name>IN_2</name></connection>
<intersection>92.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-47.5,100,-47.5</points>
<connection>
<GID>57</GID>
<name>OUT_1</name></connection>
<intersection>87.5 31</intersection>
<intersection>100 25</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>100,-47.5,100,-26</points>
<intersection>-47.5 1</intersection>
<intersection>-34 30</intersection>
<intersection>-26 26</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>100,-26,108,-26</points>
<connection>
<GID>61</GID>
<name>IN_B_2</name></connection>
<intersection>100 25</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>100,-34,108,-34</points>
<connection>
<GID>61</GID>
<name>IN_3</name></connection>
<intersection>100 25</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>87.5,-55,87.5,-47.5</points>
<intersection>-55 32</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>87.5,-55,94.5,-55</points>
<connection>
<GID>251</GID>
<name>IN_1</name></connection>
<intersection>87.5 31</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-21,111,-21</points>
<connection>
<GID>61</GID>
<name>carry_in</name></connection>
<connection>
<GID>60</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-37,111,-37</points>
<connection>
<GID>61</GID>
<name>carry_out</name></connection>
<connection>
<GID>62</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-12.5,135.5,-11.5</points>
<intersection>-12.5 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-12.5,155.5,-12.5</points>
<connection>
<GID>147</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-11.5,135.5,-11.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-15.5,135.5,-12.5</points>
<intersection>-15.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-15.5,155.5,-15.5</points>
<connection>
<GID>148</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-12.5,135.5,-12.5</points>
<connection>
<GID>60</GID>
<name>OUT_1</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-18.5,135.5,-13.5</points>
<intersection>-18.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-18.5,155.5,-18.5</points>
<connection>
<GID>149</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-13.5,135.5,-13.5</points>
<connection>
<GID>60</GID>
<name>OUT_2</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-21.5,135.5,-14.5</points>
<intersection>-21.5 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-21.5,155.5,-21.5</points>
<connection>
<GID>150</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-14.5,135.5,-14.5</points>
<connection>
<GID>60</GID>
<name>OUT_3</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-27.5,135.5,-26.5</points>
<intersection>-27.5 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-26.5,155.5,-26.5</points>
<connection>
<GID>151</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-27.5,135.5,-27.5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-29.5,135.5,-28.5</points>
<intersection>-29.5 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-29.5,155.5,-29.5</points>
<connection>
<GID>152</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-28.5,135.5,-28.5</points>
<connection>
<GID>61</GID>
<name>OUT_1</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-32.5,135.5,-29.5</points>
<intersection>-32.5 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-32.5,155.5,-32.5</points>
<connection>
<GID>153</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-29.5,135.5,-29.5</points>
<connection>
<GID>61</GID>
<name>OUT_2</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-35.5,135.5,-30.5</points>
<intersection>-35.5 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-35.5,155.5,-35.5</points>
<connection>
<GID>154</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-30.5,135.5,-30.5</points>
<connection>
<GID>61</GID>
<name>OUT_3</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-43.5,135.5,-39.5</points>
<intersection>-43.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-39.5,155.5,-39.5</points>
<connection>
<GID>155</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-43.5,135.5,-43.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-44.5,135.5,-42.5</points>
<intersection>-44.5 2</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-42.5,155.5,-42.5</points>
<connection>
<GID>156</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-44.5,135.5,-44.5</points>
<connection>
<GID>62</GID>
<name>OUT_1</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-45.5,155.5,-45.5</points>
<connection>
<GID>157</GID>
<name>N_in0</name></connection>
<connection>
<GID>62</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-48.5,135.5,-46.5</points>
<intersection>-48.5 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-48.5,155.5,-48.5</points>
<connection>
<GID>158</GID>
<name>N_in0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-46.5,135.5,-46.5</points>
<connection>
<GID>62</GID>
<name>OUT_3</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-46.5,95,-25</points>
<intersection>-46.5 2</intersection>
<intersection>-33 4</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-25,108,-25</points>
<connection>
<GID>61</GID>
<name>IN_B_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-46.5,95,-46.5</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>91.5 5</intersection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>95,-33,108,-33</points>
<connection>
<GID>61</GID>
<name>IN_2</name></connection>
<intersection>95 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>91.5,-56,91.5,-46.5</points>
<intersection>-56 6</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>91.5,-56,94.5,-56</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>91.5 5</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 2>
<page 3>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 3>
<page 4>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 4>
<page 5>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 5>
<page 6>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 6>
<page 7>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 7>
<page 8>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 8>
<page 9>
<PageViewport>0,232.907,1778,-694.093</PageViewport></page 9></circuit>