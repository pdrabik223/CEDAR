<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-46.186,-47.6584,75.6827,-184.761</PageViewport>
<gate>
<ID>2</ID>
<type>BE_NOR2</type>
<position>17.5,-9.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>-0.5,-8</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>-0.5,-17.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>GA_LED</type>
<position>23.5,-16</position>
<input>
<ID>N_in0</ID>6 </input>
<input>
<ID>N_in1</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>23.5,-19.5</position>
<input>
<ID>N_in0</ID>10 </input>
<input>
<ID>N_in1</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>GA_LED</type>
<position>25.5,-9.5</position>
<input>
<ID>N_in0</ID>12 </input>
<input>
<ID>N_in1</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>BA_NAND2</type>
<position>30,-17</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>25.5,-6</position>
<gparam>LABEL_TEXT U</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AE_SMALL_INVERTER</type>
<position>18.5,-18</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_SMALL_INVERTER</type>
<position>18.5,-16</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>31,-9.5</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>23.5,-13</position>
<gparam>LABEL_TEXT V</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>5.5,-8.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>23.5,-21.5</position>
<gparam>LABEL_TEXT W</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>5.5,-18</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>36.5,-16.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>34,-9.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>36.5,-9</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>34,-17</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>3,-55</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>19,-3</position>
<gparam>LABEL_TEXT zadanie 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>3,-64.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>15.5,-55.5</position>
<input>
<ID>N_in0</ID>15 </input>
<input>
<ID>N_in1</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>15.5,-52.5</position>
<gparam>LABEL_TEXT !A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>26,-56.5</position>
<input>
<ID>N_in0</ID>17 </input>
<input>
<ID>N_in1</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>26,-58.5</position>
<gparam>LABEL_TEXT W</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>38.5,-63.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>38.5,-56</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>39.5,-86</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>39.5,-78.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>4,-78</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>4,-87.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>23,-86</position>
<input>
<ID>N_in0</ID>21 </input>
<input>
<ID>N_in1</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>23,-89.5</position>
<input>
<ID>N_in0</ID>22 </input>
<input>
<ID>N_in1</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>25,-79.5</position>
<input>
<ID>N_in0</ID>20 </input>
<input>
<ID>N_in1</ID>18 </input>
<input>
<ID>N_in2</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>25,-76</position>
<gparam>LABEL_TEXT U</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>23,-83</position>
<gparam>LABEL_TEXT V</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>23,-91.5</position>
<gparam>LABEL_TEXT W</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>4,-127.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>4,-131</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>7,-55.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>7,-65</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>35.5,-56.5</position>
<input>
<ID>N_in0</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>GA_LED</type>
<position>35.5,-64</position>
<input>
<ID>N_in0</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>20.5,-48</position>
<gparam>LABEL_TEXT zadanie 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>4,-134.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>51,-143.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>50,-131.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>34.5,-141.5</position>
<input>
<ID>N_in0</ID>25 </input>
<input>
<ID>N_in1</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>32.5,-134</position>
<input>
<ID>N_in0</ID>27 </input>
<input>
<ID>N_in1</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>32.5,-129</position>
<input>
<ID>N_in0</ID>30 </input>
<input>
<ID>N_in1</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AE_SMALL_INVERTER</type>
<position>11,-55.5</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>32.5,-126</position>
<gparam>LABEL_TEXT U</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>BE_NOR2</type>
<position>21,-56.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AE_SMALL_INVERTER</type>
<position>30.5,-56.5</position>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>57</ID>
<type>AE_SMALL_INVERTER</type>
<position>18.5,-65</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>32.5,-136</position>
<gparam>LABEL_TEXT V</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>BA_NAND2</type>
<position>31.5,-64</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>8,-78.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_TOGGLE</type>
<position>8,-88</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>36.5,-79.5</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>GA_LED</type>
<position>36.5,-87</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>21.5,-71.5</position>
<gparam>LABEL_TEXT zadanie 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>35,-138.5</position>
<gparam>LABEL_TEXT W</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>BA_NAND2</type>
<position>17.5,-79.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_SMALL_INVERTER</type>
<position>32,-79.5</position>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_SMALL_INVERTER</type>
<position>17,-86</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_SMALL_INVERTER</type>
<position>17,-88</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>74</ID>
<type>BE_NOR2</type>
<position>30.5,-87</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>22.5,-122</position>
<gparam>LABEL_TEXT zadanie 5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>7,-128</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_TOGGLE</type>
<position>7,-131.5</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>7,-135</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>96</ID>
<type>BA_NAND2</type>
<position>24.5,-129</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_SMALL_INVERTER</type>
<position>29.5,-129</position>
<input>
<ID>IN_0</ID>53 </input>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>98</ID>
<type>BA_NAND2</type>
<position>24.5,-134</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_SMALL_INVERTER</type>
<position>29.5,-134</position>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>101</ID>
<type>BE_NOR2</type>
<position>38.5,-132</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_SMALL_INVERTER</type>
<position>43.5,-132</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>103</ID>
<type>GA_LED</type>
<position>46.5,-132</position>
<input>
<ID>N_in0</ID>58 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AE_SMALL_INVERTER</type>
<position>23.5,-140</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AE_SMALL_INVERTER</type>
<position>23.5,-143</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>106</ID>
<type>BA_NAND2</type>
<position>30.5,-141.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>BA_NAND2</type>
<position>39,-144</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AE_SMALL_INVERTER</type>
<position>44,-144</position>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>109</ID>
<type>GA_LED</type>
<position>48,-144</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-19.5,27,-19.5</points>
<connection>
<GID>6</GID>
<name>N_in1</name></connection>
<intersection>27 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>27,-19.5,27,-18</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>-19.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-16,27,-16</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-16,22.5,-16</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<connection>
<GID>5</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-18,16.5,-18</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>14.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14.5,-18,14.5,-10.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-18 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>33,-9.5,33,-9.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>18</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>33,-17,33,-17</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-19.5,22.5,-19.5</points>
<connection>
<GID>6</GID>
<name>N_in0</name></connection>
<intersection>20.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>20.5,-19.5,20.5,-18</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-9.5,29,-9.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>7</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-9.5,24.5,-9.5</points>
<connection>
<GID>7</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-55.5,18,-55.5</points>
<connection>
<GID>24</GID>
<name>N_in1</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-55.5,14.5,-55.5</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-56.5,28.5,-56.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-56.5,25,-56.5</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<connection>
<GID>55</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-79.5,30,-79.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>N_in1</name></connection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-80.5,25,-79.5</points>
<connection>
<GID>36</GID>
<name>N_in2</name></connection>
<intersection>-79.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-8.5,14.5,-8.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>12 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>12,-16,12,-8.5</points>
<intersection>-16 4</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>12,-16,16.5,-16</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>12 3</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-79.5,24,-79.5</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<connection>
<GID>36</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-86,22,-86</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<connection>
<GID>34</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-89.5,20.5,-88</points>
<intersection>-89.5 1</intersection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-89.5,22,-89.5</points>
<connection>
<GID>35</GID>
<name>N_in0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-88,20.5,-88</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-89.5,25.5,-88</points>
<intersection>-89.5 2</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-88,27.5,-88</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-89.5,25.5,-89.5</points>
<connection>
<GID>35</GID>
<name>N_in1</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-86,27.5,-86</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-141.5,33.5,-141.5</points>
<connection>
<GID>50</GID>
<name>N_in0</name></connection>
<connection>
<GID>106</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-143,35.5,-141.5</points>
<connection>
<GID>50</GID>
<name>N_in1</name></connection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-143,36,-143</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-134,31.5,-134</points>
<connection>
<GID>51</GID>
<name>N_in0</name></connection>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-134,34.5,-133</points>
<intersection>-134 1</intersection>
<intersection>-133 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-134,34.5,-134</points>
<connection>
<GID>51</GID>
<name>N_in1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-133,35.5,-133</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-63,9,-55.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-63,28.5,-63</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-129,31.5,-129</points>
<connection>
<GID>52</GID>
<name>N_in0</name></connection>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32.5,-56.5,34.5,-56.5</points>
<connection>
<GID>44</GID>
<name>N_in0</name></connection>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-64,34.5,-64</points>
<connection>
<GID>45</GID>
<name>N_in0</name></connection>
<connection>
<GID>59</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-65,11,-57.5</points>
<intersection>-65 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-65,16.5,-65</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-57.5,18,-57.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-65,28.5,-65</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-131,34.5,-129</points>
<intersection>-131 2</intersection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-129,34.5,-129</points>
<connection>
<GID>52</GID>
<name>N_in1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-131,35.5,-131</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-79.5,35.5,-79.5</points>
<connection>
<GID>62</GID>
<name>N_in0</name></connection>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-87,35.5,-87</points>
<connection>
<GID>63</GID>
<name>N_in0</name></connection>
<connection>
<GID>74</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-86,11.5,-78.5</points>
<intersection>-86 2</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-78.5,14.5,-78.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-86,15,-86</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-88,12.5,-80.5</points>
<intersection>-88 1</intersection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-88,15,-88</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-80.5,14.5,-80.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-129,27.5,-129</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<connection>
<GID>97</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-134,27.5,-134</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-132,41.5,-132</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-132,45.5,-132</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<connection>
<GID>103</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-140.5,26.5,-140</points>
<intersection>-140.5 2</intersection>
<intersection>-140 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-140,26.5,-140</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-140.5,27.5,-140.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-143,26.5,-142.5</points>
<intersection>-143 2</intersection>
<intersection>-142.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-142.5,27.5,-142.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-143,26.5,-143</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-144,42,-144</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-144,47,-144</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<connection>
<GID>109</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-145,10.5,-130</points>
<intersection>-145 1</intersection>
<intersection>-135 2</intersection>
<intersection>-130 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-145,36,-145</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9,-135,21.5,-135</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>10.5,-130,21.5,-130</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-143,12.5,-131.5</points>
<intersection>-143 2</intersection>
<intersection>-133 3</intersection>
<intersection>-131.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-131.5,12.5,-131.5</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-143,21.5,-143</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>12.5,-133,21.5,-133</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9,-128,21.5,-128</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>14.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>14.5,-140,14.5,-128</points>
<intersection>-140 5</intersection>
<intersection>-128 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>14.5,-140,21.5,-140</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>14.5 4</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-3.20825,0,159.284,-182.803</PageViewport></page 1>
<page 2>
<PageViewport>-3.20825,0,159.284,-182.803</PageViewport></page 2>
<page 3>
<PageViewport>-3.20825,0,159.284,-182.803</PageViewport></page 3>
<page 4>
<PageViewport>-3.20825,0,159.284,-182.803</PageViewport></page 4>
<page 5>
<PageViewport>-3.20825,0,159.284,-182.803</PageViewport></page 5>
<page 6>
<PageViewport>-3.20825,0,159.284,-182.803</PageViewport></page 6>
<page 7>
<PageViewport>-3.20825,0,159.284,-182.803</PageViewport></page 7>
<page 8>
<PageViewport>-3.20825,0,159.284,-182.803</PageViewport></page 8>
<page 9>
<PageViewport>-3.20825,0,159.284,-182.803</PageViewport></page 9></circuit>