<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>24.6333,-8.04087,447.541,-228.533</PageViewport>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>84.5,-22.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_DFF_LOW</type>
<position>127,-24</position>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>32</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>65,-15</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>34</ID>
<type>BE_JKFF_LOW</type>
<position>103.5,-35</position>
<input>
<ID>J</ID>5 </input>
<input>
<ID>K</ID>5 </input>
<output>
<ID>Q</ID>24 </output>
<input>
<ID>clock</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>46</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>58.5,-15</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>47</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>52,-15</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>56</ID>
<type>GA_LED</type>
<position>36.5,-14.5</position>
<input>
<ID>N_in0</ID>23 </input>
<input>
<ID>N_in1</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>GA_LED</type>
<position>38.5,-14.5</position>
<input>
<ID>N_in0</ID>22 </input>
<input>
<ID>N_in1</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>40.5,-14.5</position>
<input>
<ID>N_in0</ID>22 </input>
<input>
<ID>N_in1</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>42.5,-14.5</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>DA_FROM</type>
<position>33.5,-14.5</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID om</lparam></gate>
<gate>
<ID>65</ID>
<type>DE_TO</type>
<position>108.5,-33</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID om</lparam></gate>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>86.5,-35,100.5,-35</points>
<connection>
<GID>34</GID>
<name>clock</name></connection>
<intersection>86.5 3</intersection>
<intersection>100.5 18</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>86.5,-35,86.5,-22.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-35 2</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>100.5,-37,100.5,-33</points>
<connection>
<GID>34</GID>
<name>J</name></connection>
<connection>
<GID>34</GID>
<name>K</name></connection>
<intersection>-35 2</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>41.5,-14.5,41.5,-14.5</points>
<connection>
<GID>58</GID>
<name>N_in1</name></connection>
<connection>
<GID>59</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-14.5,39.5,-14.5</points>
<connection>
<GID>56</GID>
<name>N_in1</name></connection>
<connection>
<GID>57</GID>
<name>N_in0</name></connection>
<connection>
<GID>57</GID>
<name>N_in1</name></connection>
<connection>
<GID>58</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-14.5,35.5,-14.5</points>
<connection>
<GID>56</GID>
<name>N_in0</name></connection>
<connection>
<GID>60</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-33,106.5,-33</points>
<connection>
<GID>34</GID>
<name>Q</name></connection>
<connection>
<GID>65</GID>
<name>IN_0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>21.1819,54.6107,303.12,-92.3839</PageViewport>
<gate>
<ID>1</ID>
<type>AE_REGISTER8</type>
<position>128.5,-27.5</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>197 </input>
<input>
<ID>IN_2</ID>196 </input>
<input>
<ID>IN_3</ID>195 </input>
<input>
<ID>IN_4</ID>194 </input>
<input>
<ID>IN_5</ID>193 </input>
<input>
<ID>IN_6</ID>192 </input>
<input>
<ID>IN_7</ID>191 </input>
<output>
<ID>OUT_0</ID>244 </output>
<output>
<ID>OUT_1</ID>245 </output>
<output>
<ID>OUT_2</ID>246 </output>
<output>
<ID>OUT_3</ID>247 </output>
<output>
<ID>OUT_4</ID>248 </output>
<output>
<ID>OUT_5</ID>249 </output>
<output>
<ID>OUT_6</ID>250 </output>
<output>
<ID>OUT_7</ID>251 </output>
<input>
<ID>clear</ID>258 </input>
<input>
<ID>clock</ID>257 </input>
<input>
<ID>load</ID>6 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>194</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>99.5,-3</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>176 </input>
<input>
<ID>IN_2</ID>177 </input>
<input>
<ID>IN_3</ID>178 </input>
<output>
<ID>OUT_0</ID>198 </output>
<output>
<ID>OUT_1</ID>197 </output>
<output>
<ID>OUT_2</ID>196 </output>
<output>
<ID>OUT_3</ID>195 </output>
<output>
<ID>carry_out</ID>120 </output>
<input>
<ID>clear</ID>254 </input>
<input>
<ID>clock</ID>232 </input>
<input>
<ID>load</ID>10 </input>
<input>
<ID>shift_enable</ID>122 </input>
<input>
<ID>shift_left</ID>181 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>2</ID>
<type>CC_PULSE</type>
<position>19.5,-14</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3</ID>
<type>DE_TO</type>
<position>19.5,-9.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>196</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>135.5,-10</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>197 </input>
<input>
<ID>IN_2</ID>196 </input>
<input>
<ID>IN_3</ID>195 </input>
<input>
<ID>IN_4</ID>194 </input>
<input>
<ID>IN_5</ID>193 </input>
<input>
<ID>IN_6</ID>192 </input>
<input>
<ID>IN_7</ID>191 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 153</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>4</ID>
<type>DA_FROM</type>
<position>122.5,-42</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>197</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>99.5,-16</position>
<output>
<ID>OUT_0</ID>194 </output>
<output>
<ID>OUT_1</ID>193 </output>
<output>
<ID>OUT_2</ID>192 </output>
<output>
<ID>OUT_3</ID>191 </output>
<input>
<ID>carry_in</ID>120 </input>
<input>
<ID>clear</ID>254 </input>
<input>
<ID>clock</ID>232 </input>
<input>
<ID>shift_enable</ID>122 </input>
<input>
<ID>shift_left</ID>229 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>70,-23.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_SMALL_INVERTER</type>
<position>74,-23.5</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>DA_FROM</type>
<position>132,-42</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>201</ID>
<type>CC_PULSE</type>
<position>19,4</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 9</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>10</ID>
<type>AE_SMALL_INVERTER</type>
<position>86,-23.5</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_SMALL_INVERTER</type>
<position>90,-23.5</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>205</ID>
<type>BB_CLOCK</type>
<position>40.5,-26</position>
<output>
<ID>CLK</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>78,-23.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_SMALL_INVERTER</type>
<position>82,-23.5</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>15</ID>
<type>CC_PULSE</type>
<position>24,-13.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>24,-9.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>100.5,-39.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>237</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>48,-19.5</position>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUT_0</ID>167 </output>
<output>
<ID>OUT_1</ID>168 </output>
<output>
<ID>OUT_2</ID>169 </output>
<output>
<ID>OUT_3</ID>170 </output>
<output>
<ID>carry_out</ID>220 </output>
<input>
<ID>clear</ID>220 </input>
<input>
<ID>clock</ID>152 </input>
<input>
<ID>load</ID>227 </input>
<input>
<ID>shift_enable</ID>160 </input>
<input>
<ID>shift_left</ID>160 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>239</ID>
<type>EE_VDD</type>
<position>43.5,-18</position>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>243</ID>
<type>AE_OR4</type>
<position>56.5,-19.5</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>168 </input>
<input>
<ID>IN_2</ID>169 </input>
<input>
<ID>IN_3</ID>170 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>247</ID>
<type>GA_LED</type>
<position>67.5,-20.5</position>
<input>
<ID>N_in0</ID>206 </input>
<input>
<ID>N_in1</ID>174 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>249</ID>
<type>DE_TO</type>
<position>70.5,-20.5</position>
<input>
<ID>IN_0</ID>174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cc</lparam></gate>
<gate>
<ID>255</ID>
<type>EE_VDD</type>
<position>101.5,3</position>
<output>
<ID>OUT_0</ID>181 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>256</ID>
<type>EE_VDD</type>
<position>102.5,-10</position>
<output>
<ID>OUT_0</ID>229 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_AND2</type>
<position>63.5,-20.5</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>218 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>269</ID>
<type>AE_SMALL_INVERTER</type>
<position>52,-26</position>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>270</ID>
<type>AE_SMALL_INVERTER</type>
<position>56,-26</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>278</ID>
<type>DA_FROM</type>
<position>99.5,13.5</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID cc</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_FULLADDER_4BIT</type>
<position>173.5,-20</position>
<input>
<ID>IN_0</ID>244 </input>
<input>
<ID>IN_1</ID>245 </input>
<input>
<ID>IN_2</ID>246 </input>
<input>
<ID>IN_3</ID>247 </input>
<input>
<ID>IN_B_0</ID>198 </input>
<input>
<ID>IN_B_1</ID>197 </input>
<input>
<ID>IN_B_2</ID>196 </input>
<input>
<ID>IN_B_3</ID>195 </input>
<output>
<ID>OUT_0</ID>186 </output>
<output>
<ID>OUT_1</ID>188 </output>
<output>
<ID>OUT_2</ID>187 </output>
<output>
<ID>OUT_3</ID>189 </output>
<output>
<ID>carry_out</ID>223 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>280</ID>
<type>DE_TO</type>
<position>19,0.5</position>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID load</lparam></gate>
<gate>
<ID>88</ID>
<type>AE_FULLADDER_4BIT</type>
<position>241.5,-7</position>
<input>
<ID>IN_1</ID>204 </input>
<input>
<ID>IN_2</ID>204 </input>
<input>
<ID>IN_B_0</ID>186 </input>
<input>
<ID>IN_B_1</ID>188 </input>
<input>
<ID>IN_B_2</ID>187 </input>
<input>
<ID>IN_B_3</ID>189 </input>
<output>
<ID>OUT_0</ID>228 </output>
<output>
<ID>OUT_1</ID>226 </output>
<output>
<ID>OUT_2</ID>225 </output>
<output>
<ID>OUT_3</ID>224 </output>
<output>
<ID>carry_out</ID>241 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>89</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>229.5,-23.5</position>
<output>
<ID>A_less_B</ID>230 </output>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_3</ID>190 </input>
<input>
<ID>IN_B_0</ID>186 </input>
<input>
<ID>IN_B_1</ID>188 </input>
<input>
<ID>IN_B_2</ID>187 </input>
<input>
<ID>IN_B_3</ID>189 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>90</ID>
<type>EE_VDD</type>
<position>219.5,-28.5</position>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>91</ID>
<type>EE_VDD</type>
<position>220,-25.5</position>
<output>
<ID>OUT_0</ID>199 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_FULLADDER_4BIT</type>
<position>146,-55.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>249 </input>
<input>
<ID>IN_2</ID>250 </input>
<input>
<ID>IN_3</ID>251 </input>
<input>
<ID>IN_B_0</ID>194 </input>
<input>
<ID>IN_B_1</ID>193 </input>
<input>
<ID>IN_B_2</ID>192 </input>
<input>
<ID>IN_B_3</ID>191 </input>
<output>
<ID>OUT_0</ID>211 </output>
<output>
<ID>OUT_1</ID>213 </output>
<output>
<ID>OUT_2</ID>212 </output>
<output>
<ID>OUT_3</ID>214 </output>
<input>
<ID>carry_in</ID>223 </input>
<output>
<ID>carry_out</ID>240 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>95</ID>
<type>AE_FULLADDER_4BIT</type>
<position>244,-44</position>
<input>
<ID>IN_1</ID>222 </input>
<input>
<ID>IN_2</ID>222 </input>
<input>
<ID>IN_B_0</ID>211 </input>
<input>
<ID>IN_B_1</ID>213 </input>
<input>
<ID>IN_B_2</ID>212 </input>
<input>
<ID>IN_B_3</ID>214 </input>
<output>
<ID>OUT_0</ID>235 </output>
<output>
<ID>OUT_1</ID>236 </output>
<output>
<ID>OUT_2</ID>237 </output>
<output>
<ID>OUT_3</ID>238 </output>
<input>
<ID>carry_in</ID>241 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>289</ID>
<type>DE_TO</type>
<position>41.5,-6</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID zdradzieckamagda</lparam></gate>
<gate>
<ID>96</ID>
<type>DA_FROM</type>
<position>45,-2</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>97</ID>
<type>DA_FROM</type>
<position>45,0</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>291</ID>
<type>AE_SMALL_INVERTER</type>
<position>78,-26</position>
<input>
<ID>IN_0</ID>218 </input>
<output>
<ID>OUT_0</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>98</ID>
<type>DA_FROM</type>
<position>45,2</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>292</ID>
<type>AE_SMALL_INVERTER</type>
<position>82,-26</position>
<input>
<ID>IN_0</ID>231 </input>
<output>
<ID>OUT_0</ID>234 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>99</ID>
<type>DA_FROM</type>
<position>45,4</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>293</ID>
<type>AE_SMALL_INVERTER</type>
<position>86,-26</position>
<input>
<ID>IN_0</ID>234 </input>
<output>
<ID>OUT_0</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>45,6</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>294</ID>
<type>AE_SMALL_INVERTER</type>
<position>90,-26</position>
<input>
<ID>IN_0</ID>233 </input>
<output>
<ID>OUT_0</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>45,8</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>45,10</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>103</ID>
<type>DA_FROM</type>
<position>45,12</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>104</ID>
<type>DA_FROM</type>
<position>45,14</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>105</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>233,-59</position>
<output>
<ID>A_less_B</ID>239 </output>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_3</ID>215 </input>
<input>
<ID>IN_B_0</ID>211 </input>
<input>
<ID>IN_B_1</ID>213 </input>
<input>
<ID>IN_B_2</ID>212 </input>
<input>
<ID>IN_B_3</ID>214 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>106</ID>
<type>EE_VDD</type>
<position>228,-64</position>
<output>
<ID>OUT_0</ID>215 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>107</ID>
<type>AE_REGISTER8</type>
<position>79.5,-2.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>109 </input>
<input>
<ID>IN_2</ID>108 </input>
<input>
<ID>IN_3</ID>107 </input>
<output>
<ID>OUT_0</ID>175 </output>
<output>
<ID>OUT_1</ID>176 </output>
<output>
<ID>OUT_2</ID>177 </output>
<output>
<ID>OUT_3</ID>178 </output>
<input>
<ID>clock</ID>227 </input>
<input>
<ID>load</ID>227 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>108</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>254.5,-7</position>
<input>
<ID>IN_0</ID>228 </input>
<input>
<ID>IN_1</ID>226 </input>
<input>
<ID>IN_2</ID>225 </input>
<input>
<ID>IN_3</ID>224 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>109</ID>
<type>AE_OR2</type>
<position>236,-29</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>223 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>256,-44.5</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>236 </input>
<input>
<ID>IN_2</ID>237 </input>
<input>
<ID>IN_3</ID>238 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_OR2</type>
<position>238.5,-70.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AI_XOR2</type>
<position>224.5,-61</position>
<input>
<ID>IN_0</ID>242 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>EE_VDD</type>
<position>220.5,-60</position>
<output>
<ID>OUT_0</ID>242 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>115</ID>
<type>AE_OR2</type>
<position>99.5,-34.5</position>
<input>
<ID>IN_0</ID>256 </input>
<input>
<ID>IN_1</ID>255 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>DA_FROM</type>
<position>98.5,-39.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>117</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-23,5</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR2</type>
<position>127.5,-37</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>258 </input>
<output>
<ID>OUT</ID>257 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>71.5,5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>78 </input>
<input>
<ID>IN_2</ID>82 </input>
<input>
<ID>IN_3</ID>81 </input>
<output>
<ID>OUT_0</ID>110 </output>
<output>
<ID>OUT_1</ID>109 </output>
<output>
<ID>OUT_2</ID>108 </output>
<output>
<ID>OUT_3</ID>107 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>134</ID>
<type>BA_DECODER_2x4</type>
<position>4,-2</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_OR8</type>
<position>60.5,-6</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>69 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>68 </input>
<input>
<ID>IN_4</ID>64 </input>
<input>
<ID>IN_5</ID>65 </input>
<input>
<ID>IN_6</ID>66 </input>
<input>
<ID>IN_7</ID>67 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>140</ID>
<type>FF_GND</type>
<position>56.5,-4.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>145</ID>
<type>AE_OR2</type>
<position>60.5,16</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_OR4</type>
<position>59.5,2</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>80 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>79 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>148</ID>
<type>AE_OR4</type>
<position>59.5,10</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>80 </input>
<input>
<ID>IN_2</ID>66 </input>
<input>
<ID>IN_3</ID>84 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>149</ID>
<type>CC_PULSE</type>
<position>32,-13.5</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>150</ID>
<type>CC_PULSE</type>
<position>36,9</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>151</ID>
<type>CC_PULSE</type>
<position>32,9</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>152</ID>
<type>CC_PULSE</type>
<position>28,9</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>153</ID>
<type>CC_PULSE</type>
<position>36,1.5</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>154</ID>
<type>CC_PULSE</type>
<position>32,1.5</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>155</ID>
<type>CC_PULSE</type>
<position>28,1.5</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>156</ID>
<type>CC_PULSE</type>
<position>36,-6</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>157</ID>
<type>CC_PULSE</type>
<position>32,-6</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>158</ID>
<type>CC_PULSE</type>
<position>28,-6</position>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>159</ID>
<type>DE_TO</type>
<position>28,13</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>160</ID>
<type>DE_TO</type>
<position>32,13</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>161</ID>
<type>DE_TO</type>
<position>36,13</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>162</ID>
<type>DE_TO</type>
<position>28,5.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>163</ID>
<type>DE_TO</type>
<position>32,5.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>164</ID>
<type>DE_TO</type>
<position>36,5.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>165</ID>
<type>DE_TO</type>
<position>28,-2</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>166</ID>
<type>DE_TO</type>
<position>32,-2</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>167</ID>
<type>DE_TO</type>
<position>36,-2</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_TO</type>
<position>32,-9.5</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>172</ID>
<type>GA_LED</type>
<position>10.5,2</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>45,-4</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>183</ID>
<type>AE_OR4</type>
<position>68.5,-6</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>78 </input>
<input>
<ID>IN_3</ID>77 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>185</ID>
<type>AE_OR2</type>
<position>75.5,-9.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-15.5,107,-8</points>
<intersection>-15.5 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-8,130.5,-8</points>
<connection>
<GID>196</GID>
<name>IN_5</name></connection>
<intersection>107 0</intersection>
<intersection>115.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-15.5,107,-15.5</points>
<connection>
<GID>197</GID>
<name>OUT_1</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115.5,-51.5,115.5,-8</points>
<intersection>-51.5 6</intersection>
<intersection>-25.5 4</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>115.5,-25.5,124.5,-25.5</points>
<connection>
<GID>1</GID>
<name>IN_5</name></connection>
<intersection>115.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>115.5,-51.5,142,-51.5</points>
<connection>
<GID>94</GID>
<name>IN_B_1</name></connection>
<intersection>115.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-14.5,107,-9</points>
<intersection>-14.5 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-9,130.5,-9</points>
<connection>
<GID>196</GID>
<name>IN_4</name></connection>
<intersection>107 0</intersection>
<intersection>114.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-14.5,107,-14.5</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114.5,-50.5,114.5,-9</points>
<intersection>-50.5 8</intersection>
<intersection>-26.5 4</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>114.5,-26.5,124.5,-26.5</points>
<connection>
<GID>1</GID>
<name>IN_4</name></connection>
<intersection>114.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>114.5,-50.5,142,-50.5</points>
<connection>
<GID>94</GID>
<name>IN_B_0</name></connection>
<intersection>114.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>19.5,-12,19.5,-11.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-10,107,-4.5</points>
<intersection>-10 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-10,130.5,-10</points>
<connection>
<GID>196</GID>
<name>IN_3</name></connection>
<intersection>107 0</intersection>
<intersection>113.5 3</intersection>
<intersection>119 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-4.5,107,-4.5</points>
<connection>
<GID>194</GID>
<name>OUT_3</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>113.5,-27.5,113.5,-10</points>
<intersection>-27.5 4</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>113.5,-27.5,124.5,-27.5</points>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>113.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>119,-18,119,-10</points>
<intersection>-18 6</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>119,-18,169.5,-18</points>
<connection>
<GID>87</GID>
<name>IN_B_3</name></connection>
<intersection>119 5</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-26,54,-26</points>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection>
<connection>
<GID>270</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-11,107,-3.5</points>
<intersection>-11 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-11,130.5,-11</points>
<connection>
<GID>196</GID>
<name>IN_2</name></connection>
<intersection>107 0</intersection>
<intersection>112 3</intersection>
<intersection>119.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-3.5,107,-3.5</points>
<connection>
<GID>194</GID>
<name>OUT_2</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>112,-28.5,112,-11</points>
<intersection>-28.5 4</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>112,-28.5,124.5,-28.5</points>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>112 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>119.5,-17,119.5,-11</points>
<intersection>-17 6</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>119.5,-17,169.5,-17</points>
<connection>
<GID>87</GID>
<name>IN_B_2</name></connection>
<intersection>119.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-23.5,72,-23.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>7</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-12,107,-2.5</points>
<intersection>-12 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-12,130.5,-12</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>107 0</intersection>
<intersection>110.5 3</intersection>
<intersection>120 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-2.5,107,-2.5</points>
<connection>
<GID>194</GID>
<name>OUT_1</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110.5,-29.5,110.5,-12</points>
<intersection>-29.5 4</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>110.5,-29.5,124.5,-29.5</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>110.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>120,-16,120,-12</points>
<intersection>-16 6</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>120,-16,169.5,-16</points>
<connection>
<GID>87</GID>
<name>IN_B_1</name></connection>
<intersection>120 5</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-13,107,-1.5</points>
<intersection>-13 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-13,130.5,-13</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection>
<intersection>109.5 3</intersection>
<intersection>121 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-1.5,107,-1.5</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>109.5,-30.5,109.5,-13</points>
<intersection>-30.5 4</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>109.5,-30.5,124.5,-30.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>109.5 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>121,-15,121,-13</points>
<intersection>-15 9</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>121,-15,169.5,-15</points>
<connection>
<GID>87</GID>
<name>IN_B_0</name></connection>
<intersection>121 8</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,-25.5,225.5,-25.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<connection>
<GID>89</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-40,122.5,-21.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-40 6</intersection>
<intersection>-21.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>122.5,-21.5,127.5,-21.5</points>
<connection>
<GID>1</GID>
<name>load</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>122.5,-40,126.5,-40</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-23.5,88,-23.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<connection>
<GID>11</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-23.5,94,4</points>
<intersection>-23.5 5</intersection>
<intersection>4 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>94,4,100.5,4</points>
<intersection>94 0</intersection>
<intersection>100.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100.5,2,100.5,4</points>
<connection>
<GID>194</GID>
<name>load</name></connection>
<intersection>4 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>92,-23.5,94,-23.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>236,-26,236,-10</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>-11 30</intersection>
<intersection>-10 31</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>236,-11,237.5,-11</points>
<connection>
<GID>88</GID>
<name>IN_2</name></connection>
<intersection>236 2</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>236,-10,237.5,-10</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>236 2</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-19.5,60.5,-19.5</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<connection>
<GID>263</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-23.5,80,-23.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>13</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-20.5,66.5,-20.5</points>
<connection>
<GID>247</GID>
<name>N_in0</name></connection>
<connection>
<GID>263</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-23.5,76,-23.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-23.5,84,-23.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-11.5,24,-11.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>150,-54,229,-54</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<connection>
<GID>105</GID>
<name>IN_B_0</name></connection>
<intersection>217 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>217,-54,217,-39</points>
<intersection>-54 1</intersection>
<intersection>-39 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>217,-39,240,-39</points>
<connection>
<GID>95</GID>
<name>IN_B_0</name></connection>
<intersection>217 6</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>150,-56,229,-56</points>
<connection>
<GID>94</GID>
<name>OUT_2</name></connection>
<connection>
<GID>105</GID>
<name>IN_B_2</name></connection>
<intersection>219 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>219,-56,219,-41</points>
<intersection>-56 1</intersection>
<intersection>-41 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>219,-41,240,-41</points>
<connection>
<GID>95</GID>
<name>IN_B_2</name></connection>
<intersection>219 6</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>150,-55,229,-55</points>
<connection>
<GID>94</GID>
<name>OUT_1</name></connection>
<connection>
<GID>105</GID>
<name>IN_B_1</name></connection>
<intersection>218 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>218,-55,218,-40</points>
<intersection>-55 1</intersection>
<intersection>-40 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>218,-40,240,-40</points>
<connection>
<GID>95</GID>
<name>IN_B_1</name></connection>
<intersection>218 8</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>150,-57,229,-57</points>
<connection>
<GID>94</GID>
<name>OUT_3</name></connection>
<connection>
<GID>105</GID>
<name>IN_B_3</name></connection>
<intersection>220.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>220.5,-57,220.5,-42</points>
<intersection>-57 1</intersection>
<intersection>-42 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>220.5,-42,240,-42</points>
<connection>
<GID>95</GID>
<name>IN_B_3</name></connection>
<intersection>220.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-64,229,-64</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<connection>
<GID>105</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-26,60.5,-21.5</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<intersection>-26 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>58,-26,76,-26</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-24.5,48,-24.5</points>
<connection>
<GID>237</GID>
<name>clear</name></connection>
<connection>
<GID>237</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>241.5,-70.5,241.5,-53.5</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>-53.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>239,-53.5,241.5,-53.5</points>
<intersection>239 10</intersection>
<intersection>241.5 2</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>239,-53.5,239,-47</points>
<intersection>-53.5 8</intersection>
<intersection>-48 12</intersection>
<intersection>-47 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>239,-47,240,-47</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>239 10</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>239,-48,240,-48</points>
<connection>
<GID>95</GID>
<name>IN_2</name></connection>
<intersection>239 10</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-47.5,145,-27.5</points>
<connection>
<GID>94</GID>
<name>carry_in</name></connection>
<intersection>-34 1</intersection>
<intersection>-27.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-34,237,-34</points>
<intersection>145 0</intersection>
<intersection>237 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>237,-34,237,-32</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>145,-27.5,172.5,-27.5</points>
<intersection>145 0</intersection>
<intersection>172.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>172.5,-28,172.5,-27.5</points>
<connection>
<GID>87</GID>
<name>carry_out</name></connection>
<intersection>-27.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247.5,-8.5,247.5,-5</points>
<intersection>-8.5 1</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245.5,-8.5,247.5,-8.5</points>
<connection>
<GID>88</GID>
<name>OUT_3</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>247.5,-5,251.5,-5</points>
<connection>
<GID>108</GID>
<name>IN_3</name></connection>
<intersection>247.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247.5,-7.5,247.5,-6</points>
<intersection>-7.5 1</intersection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245.5,-7.5,247.5,-7.5</points>
<connection>
<GID>88</GID>
<name>OUT_2</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>247.5,-6,251.5,-6</points>
<connection>
<GID>108</GID>
<name>IN_2</name></connection>
<intersection>247.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245.5,-7,251.5,-7</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>245.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245.5,-7,245.5,-6.5</points>
<connection>
<GID>88</GID>
<name>OUT_1</name></connection>
<intersection>-7 1</intersection></vsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-14.5,49,-11.5</points>
<connection>
<GID>237</GID>
<name>load</name></connection>
<intersection>-12 1</intersection>
<intersection>-11.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-12,87,-12</points>
<intersection>49 0</intersection>
<intersection>87 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>87,-12,87,8</points>
<intersection>-12 1</intersection>
<intersection>-9.5 5</intersection>
<intersection>8 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>41.5,-11.5,49,-11.5</points>
<intersection>41.5 11</intersection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>78.5,8,87,8</points>
<intersection>78.5 7</intersection>
<intersection>87 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>78.5,-9.5,87,-9.5</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>78.5 8</intersection>
<intersection>87 2</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>78.5,3.5,78.5,8</points>
<connection>
<GID>107</GID>
<name>load</name></connection>
<intersection>8 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>78.5,-9.5,78.5,-7.5</points>
<connection>
<GID>107</GID>
<name>clock</name></connection>
<intersection>-9.5 5</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>41.5,-11.5,41.5,-8</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>-11.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248.5,-8,248.5,-5.5</points>
<intersection>-8 2</intersection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245.5,-5.5,248.5,-5.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<intersection>248.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>248.5,-8,251.5,-8</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>248.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-11,101.5,-10</points>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<connection>
<GID>197</GID>
<name>shift_left</name></connection></vsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>231.5,-32,235,-32</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>231.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>231.5,-32,231.5,-31.5</points>
<connection>
<GID>89</GID>
<name>A_less_B</name></connection>
<intersection>-32 2</intersection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-26,80,-26</points>
<connection>
<GID>291</GID>
<name>OUT_0</name></connection>
<connection>
<GID>292</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-26,104,-8</points>
<intersection>-26 8</intersection>
<intersection>-21 5</intersection>
<intersection>-8 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>100.5,-21,104,-21</points>
<connection>
<GID>197</GID>
<name>clock</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>100.5,-8,104,-8</points>
<connection>
<GID>194</GID>
<name>clock</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>92,-26,104,-26</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-26,88,-26</points>
<connection>
<GID>293</GID>
<name>OUT_0</name></connection>
<connection>
<GID>294</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-26,84,-26</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<connection>
<GID>293</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-45.5,250.5,-42.5</points>
<intersection>-45.5 2</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,-42.5,250.5,-42.5</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>250.5,-45.5,253,-45.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-44.5,250.5,-43.5</points>
<intersection>-44.5 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-44.5,253,-44.5</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>248,-43.5,250.5,-43.5</points>
<connection>
<GID>95</GID>
<name>OUT_1</name></connection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-44.5,250.5,-43.5</points>
<intersection>-44.5 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,-44.5,250.5,-44.5</points>
<connection>
<GID>95</GID>
<name>OUT_2</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>250.5,-43.5,253,-43.5</points>
<connection>
<GID>110</GID>
<name>IN_2</name></connection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-45.5,250.5,-42.5</points>
<intersection>-45.5 1</intersection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,-45.5,250.5,-45.5</points>
<connection>
<GID>95</GID>
<name>OUT_3</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>250.5,-42.5,253,-42.5</points>
<connection>
<GID>110</GID>
<name>IN_3</name></connection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,-69.5,235,-67</points>
<connection>
<GID>105</GID>
<name>A_less_B</name></connection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,-69.5,235.5,-69.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-71.5,145,-63.5</points>
<connection>
<GID>94</GID>
<name>carry_out</name></connection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-71.5,235.5,-71.5</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240.5,-36,240.5,-15</points>
<connection>
<GID>88</GID>
<name>carry_out</name></connection>
<intersection>-36 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216.5,-36,243,-36</points>
<connection>
<GID>95</GID>
<name>carry_in</name></connection>
<intersection>216.5 6</intersection>
<intersection>240.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>216.5,-62,216.5,-36</points>
<intersection>-62 7</intersection>
<intersection>-36 3</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>216.5,-62,221.5,-62</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>216.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221.5,-60,221.5,-60</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>227.5,-61,229,-61</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-30.5,141.5,-22</points>
<intersection>-30.5 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-22,169.5,-22</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-30.5,141.5,-30.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-29.5,142,-23</points>
<intersection>-29.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-23,169.5,-23</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-29.5,142,-29.5</points>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-28.5,142.5,-24</points>
<intersection>-28.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142.5,-24,169.5,-24</points>
<connection>
<GID>87</GID>
<name>IN_2</name></connection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-28.5,142.5,-28.5</points>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<intersection>142.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-27.5,143,-25</points>
<intersection>-27.5 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-27.5,143,-27.5</points>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143,-25,169.5,-25</points>
<connection>
<GID>87</GID>
<name>IN_3</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-57.5,138,-26.5</points>
<intersection>-57.5 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-26.5,138,-26.5</points>
<connection>
<GID>1</GID>
<name>OUT_4</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-57.5,142,-57.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-58.5,138.5,-25.5</points>
<intersection>-58.5 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-25.5,138.5,-25.5</points>
<connection>
<GID>1</GID>
<name>OUT_5</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,-58.5,142,-58.5</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-59.5,139,-24.5</points>
<intersection>-59.5 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-24.5,139,-24.5</points>
<connection>
<GID>1</GID>
<name>OUT_6</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139,-59.5,142,-59.5</points>
<connection>
<GID>94</GID>
<name>IN_2</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-60.5,139.5,-23.5</points>
<intersection>-60.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-23.5,139.5,-23.5</points>
<connection>
<GID>1</GID>
<name>OUT_7</name></connection>
<intersection>139.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139.5,-60.5,142,-60.5</points>
<connection>
<GID>94</GID>
<name>IN_3</name></connection>
<intersection>139.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-31.5,93,-8</points>
<intersection>-31.5 4</intersection>
<intersection>-8 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>93,-8,99.5,-8</points>
<connection>
<GID>194</GID>
<name>clear</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>93,-31.5,99.5,-31.5</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>93 0</intersection>
<intersection>99.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>99.5,-31.5,99.5,-21</points>
<connection>
<GID>197</GID>
<name>clear</name></connection>
<intersection>-31.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>100.5,-37.5,100.5,-37.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>98.5,-37.5,98.5,-37.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-34,127.5,-32.5</points>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<connection>
<GID>118</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-9.5,51,-2</points>
<intersection>-9.5 2</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-2,51,-2</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-9.5,57.5,-9.5</points>
<connection>
<GID>138</GID>
<name>IN_4</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-40,132,-32.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-40 5</intersection>
<intersection>-32.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>129.5,-32.5,132,-32.5</points>
<connection>
<GID>1</GID>
<name>clear</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>128.5,-40,132,-40</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-8.5,51.5,2</points>
<intersection>-8.5 2</intersection>
<intersection>1 3</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,2,51.5,2</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-8.5,57.5,-8.5</points>
<connection>
<GID>138</GID>
<name>IN_5</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51.5,1,56.5,1</points>
<connection>
<GID>147</GID>
<name>IN_2</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-7.5,52,9</points>
<intersection>-7.5 2</intersection>
<intersection>6 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,6,52,6</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-7.5,57.5,-7.5</points>
<connection>
<GID>138</GID>
<name>IN_6</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52,9,56.5,9</points>
<connection>
<GID>148</GID>
<name>IN_2</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-6.5,52.5,13</points>
<intersection>-6.5 2</intersection>
<intersection>5 3</intersection>
<intersection>10 1</intersection>
<intersection>13 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,10,52.5,10</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-6.5,57.5,-6.5</points>
<connection>
<GID>138</GID>
<name>IN_7</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52.5,5,56.5,5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,13,56.5,13</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-5.5,53,17</points>
<intersection>-5.5 2</intersection>
<intersection>14 1</intersection>
<intersection>17 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,14,53,14</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-5.5,57.5,-5.5</points>
<connection>
<GID>138</GID>
<name>IN_3</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>53,17,57.5,17</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-4.5,57.5,-2.5</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<connection>
<GID>138</GID>
<name>IN_2</name></connection>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-9,64.5,4</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>-9 6</intersection>
<intersection>4 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>64.5,4,68.5,4</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>64.5,-9,65.5,-9</points>
<connection>
<GID>183</GID>
<name>IN_3</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-7,64,5</points>
<intersection>-7 3</intersection>
<intersection>2 2</intersection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,5,68.5,5</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,2,64,2</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,-7,65.5,-7</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-1,51.5,0</points>
<intersection>-1 2</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,0,51.5,0</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-1,56.5,-1</points>
<connection>
<GID>147</GID>
<name>IN_3</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,3,51.5,11</points>
<intersection>3 2</intersection>
<intersection>8 1</intersection>
<intersection>11 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,8,51.5,8</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,3,56.5,3</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51.5,11,56.5,11</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,7,64.5,16</points>
<intersection>7 3</intersection>
<intersection>16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63.5,16,64.5,16</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64.5,7,68.5,7</points>
<connection>
<GID>119</GID>
<name>IN_3</name></connection>
<intersection>64.5 0</intersection>
<intersection>65.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>65.5,-3,65.5,7</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>7 3</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,6,64,10</points>
<intersection>6 1</intersection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,6,68.5,6</points>
<connection>
<GID>119</GID>
<name>IN_2</name></connection>
<intersection>64 0</intersection>
<intersection>65 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,10,64,10</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>64 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>65,-5,65,6</points>
<intersection>-5 6</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>65,-5,65.5,-5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>65 5</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,12,52,15</points>
<intersection>12 1</intersection>
<intersection>15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,12,52,12</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,15,57.5,15</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,4,51.5,7</points>
<intersection>4 1</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,4,51.5,4</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,7,56.5,7</points>
<connection>
<GID>148</GID>
<name>IN_3</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,11,28,11</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<connection>
<GID>159</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,11,32,11</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<connection>
<GID>160</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,11,36,11</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<connection>
<GID>161</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,3.5,28,3.5</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,3.5,32,3.5</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<connection>
<GID>163</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>36,3.5,36,3.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<connection>
<GID>164</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-4,28,-4</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<connection>
<GID>165</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-4,32,-4</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<connection>
<GID>166</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-4,36,-4</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<connection>
<GID>167</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-11.5,32,-11.5</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<connection>
<GID>168</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>72.5,-8.5,72.5,-6</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<connection>
<GID>185</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-10.5,50.5,-4</points>
<intersection>-10.5 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-4,50.5,-4</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-10.5,72.5,-10.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-2.5,70,1</points>
<connection>
<GID>119</GID>
<name>OUT_3</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-2.5,75.5,-2.5</points>
<connection>
<GID>107</GID>
<name>IN_3</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-3.5,71,1</points>
<connection>
<GID>119</GID>
<name>OUT_2</name></connection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-3.5,75.5,-3.5</points>
<connection>
<GID>107</GID>
<name>IN_2</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-4.5,72,1</points>
<connection>
<GID>119</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-4.5,75.5,-4.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-5.5,73,1</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-5.5,75.5,-5.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>20</ID>
<points>98,-11,98,-8</points>
<connection>
<GID>197</GID>
<name>carry_in</name></connection>
<connection>
<GID>194</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>108.5,-10.5,108.5,11.5</points>
<intersection>-10.5 20</intersection>
<intersection>11.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>99.5,11.5,108.5,11.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>99.5 22</intersection>
<intersection>108.5 1</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>99.5,-10.5,108.5,-10.5</points>
<intersection>99.5 21</intersection>
<intersection>108.5 1</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>99.5,-11,99.5,-10.5</points>
<connection>
<GID>197</GID>
<name>shift_enable</name></connection>
<intersection>-10.5 20</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>99.5,2,99.5,11.5</points>
<connection>
<GID>194</GID>
<name>shift_enable</name></connection>
<intersection>11.5 18</intersection></vsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>18</ID>
<points>49,-26,49,-24.5</points>
<connection>
<GID>237</GID>
<name>clock</name></connection>
<intersection>-26 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>44.5,-26,50,-26</points>
<connection>
<GID>205</GID>
<name>CLK</name></connection>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>49 18</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-18,44.5,-13.5</points>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>44.5,-13.5,50,-13.5</points>
<intersection>44.5 0</intersection>
<intersection>48 14</intersection>
<intersection>50 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>50,-14.5,50,-13.5</points>
<connection>
<GID>237</GID>
<name>shift_left</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>48,-14.5,48,-13.5</points>
<connection>
<GID>237</GID>
<name>shift_enable</name></connection>
<intersection>-13.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-18,52,-16.5</points>
<intersection>-18 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-18,52,-18</points>
<connection>
<GID>237</GID>
<name>OUT_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-16.5,53.5,-16.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-19,53.5,-19</points>
<connection>
<GID>237</GID>
<name>OUT_1</name></connection>
<intersection>53.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>53.5,-19,53.5,-18.5</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>-19 1</intersection></vsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-20.5,53.5,-20.5</points>
<connection>
<GID>243</GID>
<name>IN_2</name></connection>
<intersection>51.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>51.5,-20.5,51.5,-20</points>
<connection>
<GID>237</GID>
<name>OUT_2</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-23.5,51.5,-21</points>
<connection>
<GID>237</GID>
<name>OUT_3</name></connection>
<intersection>-23.5 12</intersection>
<intersection>-22.5 15</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>51.5,-23.5,68,-23.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>51.5,-22.5,53.5,-22.5</points>
<connection>
<GID>243</GID>
<name>IN_3</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-20.5,68.5,-20.5</points>
<connection>
<GID>247</GID>
<name>N_in1</name></connection>
<connection>
<GID>249</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-5.5,89.5,-1.5</points>
<intersection>-5.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-5.5,89.5,-5.5</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-1.5,96,-1.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-4.5,89.5,-2.5</points>
<intersection>-4.5 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-4.5,89.5,-4.5</points>
<connection>
<GID>107</GID>
<name>OUT_1</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-2.5,96,-2.5</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-3.5,96,-3.5</points>
<connection>
<GID>107</GID>
<name>OUT_2</name></connection>
<connection>
<GID>194</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-4.5,89.5,-2.5</points>
<intersection>-4.5 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-2.5,89.5,-2.5</points>
<connection>
<GID>107</GID>
<name>OUT_3</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-4.5,96,-4.5</points>
<connection>
<GID>194</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,2,101.5,2</points>
<connection>
<GID>194</GID>
<name>shift_left</name></connection>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177.5,-18.5,225.5,-18.5</points>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<connection>
<GID>89</GID>
<name>IN_B_0</name></connection>
<intersection>214.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>214.5,-18.5,214.5,-2</points>
<intersection>-18.5 1</intersection>
<intersection>-2 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>214.5,-2,237.5,-2</points>
<connection>
<GID>88</GID>
<name>IN_B_0</name></connection>
<intersection>214.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177.5,-20.5,225.5,-20.5</points>
<connection>
<GID>87</GID>
<name>OUT_2</name></connection>
<connection>
<GID>89</GID>
<name>IN_B_2</name></connection>
<intersection>216.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>216.5,-20.5,216.5,-4</points>
<intersection>-20.5 1</intersection>
<intersection>-4 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>216.5,-4,237.5,-4</points>
<connection>
<GID>88</GID>
<name>IN_B_2</name></connection>
<intersection>216.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177.5,-19.5,225.5,-19.5</points>
<connection>
<GID>87</GID>
<name>OUT_1</name></connection>
<connection>
<GID>89</GID>
<name>IN_B_1</name></connection>
<intersection>215.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>215.5,-19.5,215.5,-3</points>
<intersection>-19.5 1</intersection>
<intersection>-3 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>215.5,-3,237.5,-3</points>
<connection>
<GID>88</GID>
<name>IN_B_1</name></connection>
<intersection>215.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177.5,-21.5,225.5,-21.5</points>
<connection>
<GID>87</GID>
<name>OUT_3</name></connection>
<connection>
<GID>89</GID>
<name>IN_B_3</name></connection>
<intersection>218 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>218,-21.5,218,-5</points>
<intersection>-21.5 1</intersection>
<intersection>-5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>218,-5,237.5,-5</points>
<connection>
<GID>88</GID>
<name>IN_B_3</name></connection>
<intersection>218 6</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220.5,-28.5,225.5,-28.5</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<connection>
<GID>89</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-17.5,107,-6</points>
<intersection>-17.5 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-6,130.5,-6</points>
<connection>
<GID>196</GID>
<name>IN_7</name></connection>
<intersection>107 0</intersection>
<intersection>118 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-17.5,107,-17.5</points>
<connection>
<GID>197</GID>
<name>OUT_3</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>118,-53.5,118,-6</points>
<intersection>-53.5 6</intersection>
<intersection>-23.5 4</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>118,-23.5,124.5,-23.5</points>
<connection>
<GID>1</GID>
<name>IN_7</name></connection>
<intersection>118 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>118,-53.5,142,-53.5</points>
<connection>
<GID>94</GID>
<name>IN_B_3</name></connection>
<intersection>118 3</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-16.5,107,-7</points>
<intersection>-16.5 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-7,130.5,-7</points>
<connection>
<GID>196</GID>
<name>IN_6</name></connection>
<intersection>107 0</intersection>
<intersection>117 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-16.5,107,-16.5</points>
<connection>
<GID>197</GID>
<name>OUT_2</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>117,-52.5,117,-7</points>
<intersection>-52.5 6</intersection>
<intersection>-24.5 4</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>117,-24.5,124.5,-24.5</points>
<connection>
<GID>1</GID>
<name>IN_6</name></connection>
<intersection>117 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>117,-52.5,142,-52.5</points>
<connection>
<GID>94</GID>
<name>IN_B_2</name></connection>
<intersection>117 3</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-45.7134,30.1132,204.899,-100.549</PageViewport>
<gate>
<ID>17</ID>
<type>DD_KEYPAD_HEX</type>
<position>52,-33.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<output>
<ID>OUT_1</ID>21 </output>
<output>
<ID>OUT_2</ID>26 </output>
<output>
<ID>OUT_3</ID>27 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>19</ID>
<type>DD_KEYPAD_HEX</type>
<position>25.5,-45.5</position>
<output>
<ID>OUT_0</ID>96 </output>
<output>
<ID>OUT_1</ID>95 </output>
<output>
<ID>OUT_2</ID>76 </output>
<output>
<ID>OUT_3</ID>75 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_FULLADDER_4BIT</type>
<position>80,-39</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>95 </input>
<input>
<ID>IN_2</ID>76 </input>
<input>
<ID>IN_3</ID>75 </input>
<input>
<ID>IN_B_0</ID>19 </input>
<input>
<ID>IN_B_1</ID>21 </input>
<input>
<ID>IN_B_2</ID>26 </input>
<input>
<ID>IN_B_3</ID>27 </input>
<output>
<ID>OUT_0</ID>59 </output>
<output>
<ID>OUT_1</ID>61 </output>
<output>
<ID>OUT_2</ID>60 </output>
<output>
<ID>OUT_3</ID>62 </output>
<output>
<ID>carry_out</ID>131 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_FULLADDER_4BIT</type>
<position>129,-26</position>
<input>
<ID>IN_1</ID>97 </input>
<input>
<ID>IN_2</ID>97 </input>
<input>
<ID>IN_B_0</ID>59 </input>
<input>
<ID>IN_B_1</ID>61 </input>
<input>
<ID>IN_B_2</ID>60 </input>
<input>
<ID>IN_B_3</ID>62 </input>
<output>
<ID>OUT_0</ID>149 </output>
<output>
<ID>OUT_1</ID>148 </output>
<output>
<ID>OUT_2</ID>147 </output>
<output>
<ID>OUT_3</ID>146 </output>
<output>
<ID>carry_out</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>37</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>117,-42.5</position>
<output>
<ID>A_less_B</ID>151 </output>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_B_0</ID>59 </input>
<input>
<ID>IN_B_1</ID>61 </input>
<input>
<ID>IN_B_2</ID>60 </input>
<input>
<ID>IN_B_3</ID>62 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>39</ID>
<type>EE_VDD</type>
<position>107,-47.5</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>EE_VDD</type>
<position>107.5,-44.5</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>51</ID>
<type>DD_KEYPAD_HEX</type>
<position>52.5,-70</position>
<output>
<ID>OUT_0</ID>104 </output>
<output>
<ID>OUT_1</ID>105 </output>
<output>
<ID>OUT_2</ID>106 </output>
<output>
<ID>OUT_3</ID>111 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>52</ID>
<type>DD_KEYPAD_HEX</type>
<position>28,-82</position>
<output>
<ID>OUT_0</ID>123 </output>
<output>
<ID>OUT_1</ID>121 </output>
<output>
<ID>OUT_2</ID>119 </output>
<output>
<ID>OUT_3</ID>118 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 4</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_FULLADDER_4BIT</type>
<position>80,-74.5</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>121 </input>
<input>
<ID>IN_2</ID>119 </input>
<input>
<ID>IN_3</ID>118 </input>
<input>
<ID>IN_B_0</ID>104 </input>
<input>
<ID>IN_B_1</ID>105 </input>
<input>
<ID>IN_B_2</ID>106 </input>
<input>
<ID>IN_B_3</ID>111 </input>
<output>
<ID>OUT_0</ID>112 </output>
<output>
<ID>OUT_1</ID>114 </output>
<output>
<ID>OUT_2</ID>113 </output>
<output>
<ID>OUT_3</ID>115 </output>
<input>
<ID>carry_in</ID>131 </input>
<output>
<ID>carry_out</ID>163 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_FULLADDER_4BIT</type>
<position>131.5,-63</position>
<input>
<ID>IN_1</ID>124 </input>
<input>
<ID>IN_2</ID>124 </input>
<input>
<ID>IN_B_0</ID>112 </input>
<input>
<ID>IN_B_1</ID>114 </input>
<input>
<ID>IN_B_2</ID>113 </input>
<input>
<ID>IN_B_3</ID>115 </input>
<output>
<ID>OUT_0</ID>157 </output>
<output>
<ID>OUT_1</ID>158 </output>
<output>
<ID>OUT_2</ID>159 </output>
<output>
<ID>OUT_3</ID>161 </output>
<input>
<ID>carry_in</ID>164 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>55</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>120.5,-78</position>
<output>
<ID>A_less_B</ID>162 </output>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_3</ID>116 </input>
<input>
<ID>IN_B_0</ID>112 </input>
<input>
<ID>IN_B_1</ID>114 </input>
<input>
<ID>IN_B_2</ID>113 </input>
<input>
<ID>IN_B_3</ID>115 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>61</ID>
<type>EE_VDD</type>
<position>115.5,-83</position>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>70</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>142,-26</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>148 </input>
<input>
<ID>IN_2</ID>147 </input>
<input>
<ID>IN_3</ID>146 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_OR2</type>
<position>123.5,-48</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>143.5,-63.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>158 </input>
<input>
<ID>IN_2</ID>159 </input>
<input>
<ID>IN_3</ID>161 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_OR2</type>
<position>126,-89.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>163 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>AI_XOR2</type>
<position>112,-80</position>
<input>
<ID>IN_0</ID>166 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>EE_VDD</type>
<position>108,-79</position>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-36.5,66.5,-34</points>
<intersection>-36.5 3</intersection>
<intersection>-34 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>57,-36.5,66.5,-36.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-34,76,-34</points>
<connection>
<GID>22</GID>
<name>IN_B_0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-35,66.5,-34.5</points>
<intersection>-35 6</intersection>
<intersection>-34.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>57,-34.5,66.5,-34.5</points>
<connection>
<GID>17</GID>
<name>OUT_1</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>66.5,-35,76,-35</points>
<connection>
<GID>22</GID>
<name>IN_B_1</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-36,66.5,-32.5</points>
<intersection>-36 4</intersection>
<intersection>-32.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>57,-32.5,66.5,-32.5</points>
<connection>
<GID>17</GID>
<name>OUT_2</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-36,76,-36</points>
<connection>
<GID>22</GID>
<name>IN_B_2</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-37,66.5,-30.5</points>
<intersection>-37 4</intersection>
<intersection>-30.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>57,-30.5,66.5,-30.5</points>
<connection>
<GID>17</GID>
<name>OUT_3</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-37,76,-37</points>
<connection>
<GID>22</GID>
<name>IN_B_3</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-37.5,113,-37.5</points>
<connection>
<GID>37</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>92.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>92.5,-37.5,92.5,-21</points>
<intersection>-37.5 1</intersection>
<intersection>-21 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>92.5,-21,125,-21</points>
<connection>
<GID>27</GID>
<name>IN_B_0</name></connection>
<intersection>92.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-39.5,113,-39.5</points>
<connection>
<GID>37</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>22</GID>
<name>OUT_2</name></connection>
<intersection>94.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>94.5,-39.5,94.5,-23</points>
<intersection>-39.5 1</intersection>
<intersection>-23 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>94.5,-23,125,-23</points>
<connection>
<GID>27</GID>
<name>IN_B_2</name></connection>
<intersection>94.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-38.5,113,-38.5</points>
<connection>
<GID>37</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>22</GID>
<name>OUT_1</name></connection>
<intersection>93.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>93.5,-38.5,93.5,-22</points>
<intersection>-38.5 1</intersection>
<intersection>-22 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>93.5,-22,125,-22</points>
<connection>
<GID>27</GID>
<name>IN_B_1</name></connection>
<intersection>93.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-40.5,113,-40.5</points>
<connection>
<GID>37</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>22</GID>
<name>OUT_3</name></connection>
<intersection>96 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>96,-40.5,96,-24</points>
<intersection>-40.5 1</intersection>
<intersection>-24 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>96,-24,125,-24</points>
<connection>
<GID>27</GID>
<name>IN_B_3</name></connection>
<intersection>96 6</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-47.5,113,-47.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108.5,-44.5,113,-44.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-44,53,-42.5</points>
<intersection>-44 4</intersection>
<intersection>-42.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-42.5,53,-42.5</points>
<connection>
<GID>19</GID>
<name>OUT_3</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>53,-44,76,-44</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-44.5,53,-43</points>
<intersection>-44.5 3</intersection>
<intersection>-43 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-44.5,53,-44.5</points>
<connection>
<GID>19</GID>
<name>OUT_2</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>53,-43,76,-43</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-46.5,53,-42</points>
<intersection>-46.5 3</intersection>
<intersection>-42 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-46.5,53,-46.5</points>
<connection>
<GID>19</GID>
<name>OUT_1</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>53,-42,76,-42</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-48.5,53,-41</points>
<intersection>-48.5 3</intersection>
<intersection>-41 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-48.5,53,-48.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>53,-41,76,-41</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>123.5,-45,123.5,-29</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>-30 30</intersection>
<intersection>-29 31</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>123.5,-30,125,-30</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>123.5 2</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>123.5,-29,125,-29</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>123.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-73,66.5,-69.5</points>
<intersection>-73 3</intersection>
<intersection>-69.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>57.5,-73,66.5,-73</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-69.5,76,-69.5</points>
<connection>
<GID>53</GID>
<name>IN_B_0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-71,66.5,-70.5</points>
<intersection>-71 7</intersection>
<intersection>-70.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>57.5,-71,66.5,-71</points>
<connection>
<GID>51</GID>
<name>OUT_1</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>66.5,-70.5,76,-70.5</points>
<connection>
<GID>53</GID>
<name>IN_B_1</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-71.5,66.5,-69</points>
<intersection>-71.5 4</intersection>
<intersection>-69 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>57.5,-69,66.5,-69</points>
<connection>
<GID>51</GID>
<name>OUT_2</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-71.5,76,-71.5</points>
<connection>
<GID>53</GID>
<name>IN_B_2</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-72.5,66.5,-67</points>
<intersection>-72.5 4</intersection>
<intersection>-67 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>57.5,-67,66.5,-67</points>
<connection>
<GID>51</GID>
<name>OUT_3</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-72.5,76,-72.5</points>
<connection>
<GID>53</GID>
<name>IN_B_3</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-73,116.5,-73</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<connection>
<GID>55</GID>
<name>IN_B_0</name></connection>
<intersection>95 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>95,-73,95,-58</points>
<intersection>-73 1</intersection>
<intersection>-58 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>95,-58,127.5,-58</points>
<connection>
<GID>54</GID>
<name>IN_B_0</name></connection>
<intersection>95 6</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-75,116.5,-75</points>
<connection>
<GID>53</GID>
<name>OUT_2</name></connection>
<connection>
<GID>55</GID>
<name>IN_B_2</name></connection>
<intersection>97 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>97,-75,97,-60</points>
<intersection>-75 1</intersection>
<intersection>-60 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>97,-60,127.5,-60</points>
<connection>
<GID>54</GID>
<name>IN_B_2</name></connection>
<intersection>97 6</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-74,116.5,-74</points>
<connection>
<GID>53</GID>
<name>OUT_1</name></connection>
<connection>
<GID>55</GID>
<name>IN_B_1</name></connection>
<intersection>96 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>96,-74,96,-59</points>
<intersection>-74 1</intersection>
<intersection>-59 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>96,-59,127.5,-59</points>
<connection>
<GID>54</GID>
<name>IN_B_1</name></connection>
<intersection>96 8</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-76,116.5,-76</points>
<connection>
<GID>53</GID>
<name>OUT_3</name></connection>
<connection>
<GID>55</GID>
<name>IN_B_3</name></connection>
<intersection>98.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>98.5,-76,98.5,-61</points>
<intersection>-76 1</intersection>
<intersection>-61 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>98.5,-61,127.5,-61</points>
<connection>
<GID>54</GID>
<name>IN_B_3</name></connection>
<intersection>98.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>116.5,-83,116.5,-83</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<connection>
<GID>55</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-79.5,54.5,-79</points>
<intersection>-79.5 5</intersection>
<intersection>-79 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33,-79,54.5,-79</points>
<connection>
<GID>52</GID>
<name>OUT_3</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54.5,-79.5,76,-79.5</points>
<connection>
<GID>53</GID>
<name>IN_3</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-81,54.5,-78.5</points>
<intersection>-81 3</intersection>
<intersection>-78.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>33,-81,54.5,-81</points>
<connection>
<GID>52</GID>
<name>OUT_2</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>54.5,-78.5,76,-78.5</points>
<connection>
<GID>53</GID>
<name>IN_2</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-83,54.5,-77.5</points>
<intersection>-83 3</intersection>
<intersection>-77.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>33,-83,54.5,-83</points>
<connection>
<GID>52</GID>
<name>OUT_1</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>54.5,-77.5,76,-77.5</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-85,54.5,-76.5</points>
<intersection>-85 3</intersection>
<intersection>-76.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>33,-85,54.5,-85</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>54.5,-76.5,76,-76.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>129,-89.5,129,-72.5</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>-72.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>126.5,-72.5,129,-72.5</points>
<intersection>126.5 10</intersection>
<intersection>129 2</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>126.5,-72.5,126.5,-66</points>
<intersection>-72.5 8</intersection>
<intersection>-67 12</intersection>
<intersection>-66 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>126.5,-66,127.5,-66</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>126.5 10</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>126.5,-67,127.5,-67</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>126.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-66.5,79,-47</points>
<connection>
<GID>22</GID>
<name>carry_out</name></connection>
<connection>
<GID>53</GID>
<name>carry_in</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-53.5,124.5,-53.5</points>
<intersection>79 0</intersection>
<intersection>124.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124.5,-53.5,124.5,-51</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>-53.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-27.5,135,-24</points>
<intersection>-27.5 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-27.5,135,-27.5</points>
<connection>
<GID>27</GID>
<name>OUT_3</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135,-24,139,-24</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-26.5,135,-25</points>
<intersection>-26.5 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-26.5,135,-26.5</points>
<connection>
<GID>27</GID>
<name>OUT_2</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135,-25,139,-25</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-26,139,-26</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>133 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>133,-26,133,-25.5</points>
<connection>
<GID>27</GID>
<name>OUT_1</name></connection>
<intersection>-26 1</intersection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-27,136,-24.5</points>
<intersection>-27 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-24.5,136,-24.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>136,-27,139,-27</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>119,-51,122.5,-51</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>119 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>119,-51,119,-50.5</points>
<connection>
<GID>37</GID>
<name>A_less_B</name></connection>
<intersection>-51 2</intersection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-64.5,138,-61.5</points>
<intersection>-64.5 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-61.5,138,-61.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-64.5,140.5,-64.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-63.5,138,-62.5</points>
<intersection>-63.5 1</intersection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-63.5,140.5,-63.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135.5,-62.5,138,-62.5</points>
<connection>
<GID>54</GID>
<name>OUT_1</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-63.5,138,-62.5</points>
<intersection>-63.5 1</intersection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-63.5,138,-63.5</points>
<connection>
<GID>54</GID>
<name>OUT_2</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-62.5,140.5,-62.5</points>
<connection>
<GID>73</GID>
<name>IN_2</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-64.5,138,-61.5</points>
<intersection>-64.5 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-64.5,138,-64.5</points>
<connection>
<GID>54</GID>
<name>OUT_3</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-61.5,140.5,-61.5</points>
<connection>
<GID>73</GID>
<name>IN_3</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-88.5,122.5,-86</points>
<connection>
<GID>55</GID>
<name>A_less_B</name></connection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-88.5,123,-88.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-90.5,79,-82.5</points>
<connection>
<GID>53</GID>
<name>carry_out</name></connection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-90.5,123,-90.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-55,128,-34</points>
<connection>
<GID>27</GID>
<name>carry_out</name></connection>
<intersection>-55 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-55,130.5,-55</points>
<connection>
<GID>54</GID>
<name>carry_in</name></connection>
<intersection>104 6</intersection>
<intersection>128 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>104,-81,104,-55</points>
<intersection>-81 7</intersection>
<intersection>-55 3</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>104,-81,109,-81</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>104 6</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-79,109,-79</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>115,-80,116.5,-80</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>78</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-3.31105e-006,0.219346,317.181,-165.15</PageViewport></page 3>
<page 4>
<PageViewport>-3.31105e-006,0.219346,317.181,-165.15</PageViewport></page 4>
<page 5>
<PageViewport>-3.31105e-006,0.219346,317.181,-165.15</PageViewport></page 5>
<page 6>
<PageViewport>-3.31105e-006,0.219346,317.181,-165.15</PageViewport></page 6>
<page 7>
<PageViewport>-3.31105e-006,0.219346,317.181,-165.15</PageViewport></page 7>
<page 8>
<PageViewport>-3.31105e-006,0.219346,317.181,-165.15</PageViewport></page 8>
<page 9>
<PageViewport>-3.31105e-006,0.219346,317.181,-165.15</PageViewport></page 9></circuit>