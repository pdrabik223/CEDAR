<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-163.383,61.7175,399.148,-231.571</PageViewport>
<gate>
<ID>2</ID>
<type>BE_NOR2</type>
<position>22.5,-31</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>4.5,-29.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>4.5,-39</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>GA_LED</type>
<position>28.5,-37.5</position>
<input>
<ID>N_in0</ID>6 </input>
<input>
<ID>N_in1</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>28.5,-41</position>
<input>
<ID>N_in0</ID>10 </input>
<input>
<ID>N_in1</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>GA_LED</type>
<position>30.5,-31</position>
<input>
<ID>N_in0</ID>12 </input>
<input>
<ID>N_in1</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>BA_NAND2</type>
<position>35,-38.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>30.5,-27.5</position>
<gparam>LABEL_TEXT U</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AE_SMALL_INVERTER</type>
<position>23.5,-39.5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_SMALL_INVERTER</type>
<position>23.5,-37.5</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>36,-31</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>28.5,-34.5</position>
<gparam>LABEL_TEXT V</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>10.5,-30</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>28.5,-43</position>
<gparam>LABEL_TEXT W</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>10.5,-39.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>41.5,-38</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>39,-31</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>41.5,-30.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>39,-38.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>3,-55</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>24,-24.5</position>
<gparam>LABEL_TEXT zadanie 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>3,-64.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>15.5,-55.5</position>
<input>
<ID>N_in0</ID>15 </input>
<input>
<ID>N_in1</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>15.5,-52.5</position>
<gparam>LABEL_TEXT !A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>26,-56.5</position>
<input>
<ID>N_in0</ID>17 </input>
<input>
<ID>N_in1</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>26,-58.5</position>
<gparam>LABEL_TEXT W</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>38.5,-63.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>38.5,-56</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>39.5,-87.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>39.5,-78.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>4,-78</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>4,-89</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>23,-87.5</position>
<input>
<ID>N_in0</ID>21 </input>
<input>
<ID>N_in1</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>23,-91</position>
<input>
<ID>N_in0</ID>22 </input>
<input>
<ID>N_in1</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>25,-79.5</position>
<input>
<ID>N_in0</ID>20 </input>
<input>
<ID>N_in1</ID>18 </input>
<input>
<ID>N_in2</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>25,-76</position>
<gparam>LABEL_TEXT U</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>23,-84.5</position>
<gparam>LABEL_TEXT V</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>23,-93</position>
<gparam>LABEL_TEXT W</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>1,-109.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>1,-113</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>7,-55.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>7,-65</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>35.5,-56.5</position>
<input>
<ID>N_in0</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>GA_LED</type>
<position>35.5,-64</position>
<input>
<ID>N_in0</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>21,-48</position>
<gparam>LABEL_TEXT zadanie 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>1,-116.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>48,-125.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>47,-113.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>31.5,-123.5</position>
<input>
<ID>N_in0</ID>25 </input>
<input>
<ID>N_in1</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>29.5,-116</position>
<input>
<ID>N_in0</ID>27 </input>
<input>
<ID>N_in1</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>29.5,-111</position>
<input>
<ID>N_in0</ID>30 </input>
<input>
<ID>N_in1</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AE_SMALL_INVERTER</type>
<position>11,-55.5</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>29.5,-108</position>
<gparam>LABEL_TEXT U</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>BE_NOR2</type>
<position>21,-56.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AE_SMALL_INVERTER</type>
<position>30.5,-56.5</position>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>57</ID>
<type>AE_SMALL_INVERTER</type>
<position>18.5,-65</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>29.5,-118</position>
<gparam>LABEL_TEXT V</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>BA_NAND2</type>
<position>31.5,-64</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>8,-78.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_TOGGLE</type>
<position>8,-89.5</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>36.5,-79.5</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>GA_LED</type>
<position>36.5,-88.5</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>21.5,-71.5</position>
<gparam>LABEL_TEXT zadanie 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>32,-120.5</position>
<gparam>LABEL_TEXT W</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>BA_NAND2</type>
<position>17.5,-79.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_SMALL_INVERTER</type>
<position>32,-79.5</position>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_SMALL_INVERTER</type>
<position>17,-87.5</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_SMALL_INVERTER</type>
<position>17,-89.5</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>74</ID>
<type>BE_NOR2</type>
<position>30.5,-88.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>19.5,-104</position>
<gparam>LABEL_TEXT zadanie 5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>4,-110</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_TOGGLE</type>
<position>4,-113.5</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>4,-117</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>96</ID>
<type>BA_NAND2</type>
<position>21.5,-111</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_SMALL_INVERTER</type>
<position>26.5,-111</position>
<input>
<ID>IN_0</ID>53 </input>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>98</ID>
<type>BA_NAND2</type>
<position>21.5,-116</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_SMALL_INVERTER</type>
<position>26.5,-116</position>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>101</ID>
<type>BE_NOR2</type>
<position>35.5,-114</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_SMALL_INVERTER</type>
<position>40.5,-114</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>103</ID>
<type>GA_LED</type>
<position>43.5,-114</position>
<input>
<ID>N_in0</ID>58 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AE_SMALL_INVERTER</type>
<position>20.5,-122</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AE_SMALL_INVERTER</type>
<position>20.5,-125</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>106</ID>
<type>BA_NAND2</type>
<position>27.5,-123.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>BA_NAND2</type>
<position>36,-126</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AE_SMALL_INVERTER</type>
<position>41,-126</position>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>109</ID>
<type>GA_LED</type>
<position>45,-126</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-41,32,-41</points>
<connection>
<GID>6</GID>
<name>N_in1</name></connection>
<intersection>32 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>32,-41,32,-39.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>-41 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-37.5,32,-37.5</points>
<connection>
<GID>5</GID>
<name>N_in1</name></connection>
<connection>
<GID>8</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-37.5,27.5,-37.5</points>
<connection>
<GID>5</GID>
<name>N_in0</name></connection>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-39.5,21.5,-39.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>19.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19.5,-39.5,19.5,-32</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-39.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>38,-31,38,-31</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>18</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>38,-38.5,38,-38.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-41,27.5,-41</points>
<connection>
<GID>6</GID>
<name>N_in0</name></connection>
<intersection>25.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>25.5,-41,25.5,-39.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-41 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-31,34,-31</points>
<connection>
<GID>7</GID>
<name>N_in1</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-31,29.5,-31</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>7</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-55.5,18,-55.5</points>
<connection>
<GID>24</GID>
<name>N_in1</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-55.5,14.5,-55.5</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-56.5,28.5,-56.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-56.5,25,-56.5</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<connection>
<GID>55</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-79.5,30,-79.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>N_in1</name></connection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-80.5,25,-79.5</points>
<connection>
<GID>36</GID>
<name>N_in2</name></connection>
<intersection>-79.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-30,19.5,-30</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>17 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>17,-37.5,17,-30</points>
<intersection>-37.5 4</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>17,-37.5,21.5,-37.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>17 3</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-79.5,24,-79.5</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<connection>
<GID>36</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-87.5,22,-87.5</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-91,20.5,-89.5</points>
<intersection>-91 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-91,22,-91</points>
<connection>
<GID>35</GID>
<name>N_in0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-89.5,20.5,-89.5</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-91,25.5,-89.5</points>
<intersection>-91 2</intersection>
<intersection>-89.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24,-91,25.5,-91</points>
<connection>
<GID>35</GID>
<name>N_in1</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25.5,-89.5,27.5,-89.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-87.5,27.5,-87.5</points>
<connection>
<GID>34</GID>
<name>N_in1</name></connection>
<connection>
<GID>74</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-123.5,30.5,-123.5</points>
<connection>
<GID>50</GID>
<name>N_in0</name></connection>
<connection>
<GID>106</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-125,32.5,-123.5</points>
<connection>
<GID>50</GID>
<name>N_in1</name></connection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-125,33,-125</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-116,28.5,-116</points>
<connection>
<GID>51</GID>
<name>N_in0</name></connection>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-116,31.5,-115</points>
<intersection>-116 1</intersection>
<intersection>-115 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-116,31.5,-116</points>
<connection>
<GID>51</GID>
<name>N_in1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-115,32.5,-115</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-63,9,-55.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-63,28.5,-63</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-111,28.5,-111</points>
<connection>
<GID>52</GID>
<name>N_in0</name></connection>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32.5,-56.5,34.5,-56.5</points>
<connection>
<GID>44</GID>
<name>N_in0</name></connection>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-64,34.5,-64</points>
<connection>
<GID>45</GID>
<name>N_in0</name></connection>
<connection>
<GID>59</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-65,11,-57.5</points>
<intersection>-65 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-65,16.5,-65</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-57.5,18,-57.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-65,28.5,-65</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-113,31.5,-111</points>
<intersection>-113 3</intersection>
<intersection>-111 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-111,31.5,-111</points>
<connection>
<GID>52</GID>
<name>N_in1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-113,32.5,-113</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-79.5,35.5,-79.5</points>
<connection>
<GID>62</GID>
<name>N_in0</name></connection>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-88.5,35.5,-88.5</points>
<connection>
<GID>63</GID>
<name>N_in0</name></connection>
<connection>
<GID>74</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-87.5,11.5,-78.5</points>
<intersection>-87.5 2</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-78.5,14.5,-78.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-87.5,15,-87.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-89.5,12.5,-80.5</points>
<intersection>-89.5 1</intersection>
<intersection>-89.5 1</intersection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-89.5,15,-89.5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-80.5,14.5,-80.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-111,24.5,-111</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<connection>
<GID>97</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-116,24.5,-116</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-114,38.5,-114</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-114,42.5,-114</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<connection>
<GID>103</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-122.5,23.5,-122</points>
<intersection>-122.5 3</intersection>
<intersection>-122 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-122,23.5,-122</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23.5,-122.5,24.5,-122.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-125,23.5,-124.5</points>
<intersection>-125 2</intersection>
<intersection>-124.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-125,23.5,-125</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23.5,-124.5,24.5,-124.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-126,39,-126</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>43,-126,44,-126</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<connection>
<GID>109</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-127,7.5,-112</points>
<intersection>-127 1</intersection>
<intersection>-117 2</intersection>
<intersection>-112 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-127,33,-127</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-117,18.5,-117</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>7.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>7.5,-112,18.5,-112</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-125,9.5,-113.5</points>
<intersection>-125 2</intersection>
<intersection>-115 3</intersection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-113.5,9.5,-113.5</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-125,18.5,-125</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>9.5,-115,18.5,-115</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-110,18.5,-110</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>11.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>11.5,-122,11.5,-110</points>
<intersection>-122 5</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>11.5,-122,18.5,-122</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>11.5 4</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-10.2571,0,701.699,-371.194</PageViewport></page 1>
<page 2>
<PageViewport>-10.2571,0,701.699,-371.194</PageViewport></page 2>
<page 3>
<PageViewport>-10.2571,0,701.699,-371.194</PageViewport></page 3>
<page 4>
<PageViewport>-10.2571,0,701.699,-371.194</PageViewport></page 4>
<page 5>
<PageViewport>-10.2571,0,701.699,-371.194</PageViewport></page 5>
<page 6>
<PageViewport>-10.2571,0,701.699,-371.194</PageViewport></page 6>
<page 7>
<PageViewport>-10.2571,0,701.699,-371.194</PageViewport></page 7>
<page 8>
<PageViewport>-10.2571,0,701.699,-371.194</PageViewport></page 8>
<page 9>
<PageViewport>-10.2571,0,701.699,-371.194</PageViewport></page 9></circuit>