<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>314.786,209.74,406.69,164.314</PageViewport>
<gate>
<ID>28</ID>
<type>BB_CLOCK</type>
<position>333,183</position>
<output>
<ID>CLK</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>29</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>341,189.5</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>18 </output>
<output>
<ID>OUT_1</ID>23 </output>
<output>
<ID>OUT_2</ID>88 </output>
<output>
<ID>OUT_3</ID>89 </output>
<output>
<ID>carry_out</ID>564 </output>
<input>
<ID>clear</ID>564 </input>
<input>
<ID>clock</ID>16 </input>
<input>
<ID>load</ID>585 </input>
<input>
<ID>shift_enable</ID>17 </input>
<input>
<ID>shift_left</ID>17 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>30</ID>
<type>EE_VDD</type>
<position>336.5,191</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_OR4</type>
<position>349.5,189.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>23 </input>
<input>
<ID>IN_2</ID>88 </input>
<input>
<ID>IN_3</ID>89 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>362.5,188.5</position>
<input>
<ID>N_in0</ID>239 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>DE_TO</type>
<position>366.5,191.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cc</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND2</type>
<position>358.5,188.5</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>240 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>502</ID>
<type>GA_LED</type>
<position>342,200.5</position>
<input>
<ID>N_in2</ID>585 </input>
<input>
<ID>N_in3</ID>581 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>AE_SMALL_INVERTER</type>
<position>345,183</position>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>152</ID>
<type>AE_SMALL_INVERTER</type>
<position>349,183</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>240 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>157</ID>
<type>CC_PULSE</type>
<position>342,205</position>
<output>
<ID>OUT_0</ID>581 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 270</gparam></gate>
<wire>
<ID>581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>342,201.5,342,203</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<connection>
<GID>502</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>342,194.5,342,199.5</points>
<connection>
<GID>29</GID>
<name>load</name></connection>
<connection>
<GID>502</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347,183,347,183</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<connection>
<GID>152</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>18</ID>
<points>342,183,342,184.5</points>
<connection>
<GID>29</GID>
<name>clock</name></connection>
<intersection>183 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>337,183,343,183</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>CLK</name></connection>
<intersection>342 18</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,191,337.5,195.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>195.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>337.5,195.5,343,195.5</points>
<intersection>337.5 0</intersection>
<intersection>341 14</intersection>
<intersection>343 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>343,194.5,343,195.5</points>
<connection>
<GID>29</GID>
<name>shift_left</name></connection>
<intersection>195.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>341,194.5,341,195.5</points>
<connection>
<GID>29</GID>
<name>shift_enable</name></connection>
<intersection>195.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>345,191,345,192.5</points>
<intersection>191 1</intersection>
<intersection>192.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344.5,191,345,191</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>345 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>345,192.5,346.5,192.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>345 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>344.5,190.5,346.5,190.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>344.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>344.5,190,344.5,190.5</points>
<connection>
<GID>29</GID>
<name>OUT_1</name></connection>
<intersection>190.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361.5,188.5,361.5,188.5</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<connection>
<GID>56</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,183,355,187.5</points>
<intersection>183 5</intersection>
<intersection>187.5 15</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>351,183,355,183</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>355,187.5,355.5,187.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>344.5,188.5,346.5,188.5</points>
<connection>
<GID>31</GID>
<name>IN_2</name></connection>
<intersection>344.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>344.5,188.5,344.5,189</points>
<connection>
<GID>29</GID>
<name>OUT_2</name></connection>
<intersection>188.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344.5,186.5,344.5,188</points>
<connection>
<GID>29</GID>
<name>OUT_3</name></connection>
<intersection>186.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>344.5,186.5,346.5,186.5</points>
<connection>
<GID>31</GID>
<name>IN_3</name></connection>
<intersection>344.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>353.5,189.5,355.5,189.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>339.5,184.5,341,184.5</points>
<connection>
<GID>29</GID>
<name>clear</name></connection>
<connection>
<GID>29</GID>
<name>carry_out</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-494.141,271.986,729.859,-333.014</PageViewport></page 1>
<page 2>
<PageViewport>243.451,350.674,1467.45,-254.326</PageViewport>
<gate>
<ID>389</ID>
<type>AI_XOR2</type>
<position>334,-63</position>
<input>
<ID>IN_0</ID>530 </input>
<input>
<ID>IN_1</ID>543 </input>
<output>
<ID>OUT</ID>532 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>390</ID>
<type>AI_XOR2</type>
<position>338,-63</position>
<input>
<ID>IN_0</ID>530 </input>
<input>
<ID>IN_1</ID>542 </input>
<output>
<ID>OUT</ID>531 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>391</ID>
<type>AE_FULLADDER_4BIT</type>
<position>327,-74</position>
<input>
<ID>IN_1</ID>530 </input>
<input>
<ID>IN_3</ID>530 </input>
<input>
<ID>IN_B_0</ID>531 </input>
<input>
<ID>IN_B_1</ID>532 </input>
<input>
<ID>IN_B_2</ID>533 </input>
<input>
<ID>IN_B_3</ID>534 </input>
<output>
<ID>OUT_0</ID>541 </output>
<output>
<ID>OUT_1</ID>540 </output>
<output>
<ID>OUT_2</ID>539 </output>
<output>
<ID>OUT_3</ID>538 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>392</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>333.5,-83.5</position>
<input>
<ID>IN_0</ID>541 </input>
<input>
<ID>IN_1</ID>540 </input>
<input>
<ID>IN_2</ID>539 </input>
<input>
<ID>IN_3</ID>538 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>393</ID>
<type>GA_LED</type>
<position>324,-82.5</position>
<input>
<ID>N_in0</ID>535 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>394</ID>
<type>GA_LED</type>
<position>322,-82.5</position>
<input>
<ID>N_in0</ID>536 </input>
<input>
<ID>N_in1</ID>535 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>395</ID>
<type>GA_LED</type>
<position>320,-82.5</position>
<input>
<ID>N_in0</ID>537 </input>
<input>
<ID>N_in1</ID>536 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>396</ID>
<type>GA_LED</type>
<position>318,-82.5</position>
<input>
<ID>N_in0</ID>530 </input>
<input>
<ID>N_in1</ID>537 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>397</ID>
<type>AE_SMALL_INVERTER</type>
<position>314.5,-54.5</position>
<input>
<ID>IN_0</ID>352 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>398</ID>
<type>AI_XOR2</type>
<position>326,-37</position>
<input>
<ID>IN_0</ID>550 </input>
<input>
<ID>IN_1</ID>547 </input>
<output>
<ID>OUT</ID>546 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>399</ID>
<type>EE_VDD</type>
<position>325,-33</position>
<output>
<ID>OUT_0</ID>547 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>400</ID>
<type>AE_OR2</type>
<position>349,-49.5</position>
<input>
<ID>IN_0</ID>549 </input>
<input>
<ID>IN_1</ID>357 </input>
<output>
<ID>OUT</ID>358 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>401</ID>
<type>DD_KEYPAD_HEX</type>
<position>470.5,5.5</position>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>402</ID>
<type>DD_KEYPAD_HEX</type>
<position>470.5,17.5</position>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>403</ID>
<type>AA_AND2</type>
<position>531,30.5</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>372 </input>
<output>
<ID>OUT</ID>374 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_FULLADDER_4BIT</type>
<position>76,-35.5</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_3</ID>260 </input>
<input>
<ID>IN_B_0</ID>259 </input>
<input>
<ID>IN_B_1</ID>217 </input>
<input>
<ID>IN_B_2</ID>124 </input>
<input>
<ID>IN_B_3</ID>97 </input>
<output>
<ID>OUT_0</ID>76 </output>
<output>
<ID>OUT_1</ID>27 </output>
<output>
<ID>OUT_2</ID>26 </output>
<output>
<ID>OUT_3</ID>75 </output>
<input>
<ID>carry_in</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>404</ID>
<type>AA_AND2</type>
<position>531,19.5</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>371 </input>
<output>
<ID>OUT</ID>380 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>405</ID>
<type>AA_AND2</type>
<position>531,14</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>370 </input>
<output>
<ID>OUT</ID>402 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_AND2</type>
<position>531,9.5</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>369 </input>
<output>
<ID>OUT</ID>408 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>DD_KEYPAD_HEX</type>
<position>52,-33.5</position>
<output>
<ID>OUT_0</ID>273 </output>
<output>
<ID>OUT_1</ID>272 </output>
<output>
<ID>OUT_2</ID>271 </output>
<output>
<ID>OUT_3</ID>270 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>407</ID>
<type>AA_AND2</type>
<position>531,0</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>368 </input>
<output>
<ID>OUT</ID>410 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>63,-7</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_AND2</type>
<position>531,-4</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>351 </input>
<output>
<ID>OUT</ID>411 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>DD_KEYPAD_HEX</type>
<position>25.5,-47</position>
<output>
<ID>OUT_0</ID>106 </output>
<output>
<ID>OUT_1</ID>111 </output>
<output>
<ID>OUT_2</ID>118 </output>
<output>
<ID>OUT_3</ID>119 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_AND2</type>
<position>531,-8</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>350 </input>
<output>
<ID>OUT</ID>412 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>410</ID>
<type>AA_AND2</type>
<position>531,-12</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>314 </input>
<output>
<ID>OUT</ID>414 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>411</ID>
<type>AE_FULLADDER_4BIT</type>
<position>549.5,25.5</position>
<input>
<ID>IN_0</ID>442 </input>
<input>
<ID>IN_1</ID>441 </input>
<input>
<ID>IN_2</ID>440 </input>
<input>
<ID>IN_3</ID>425 </input>
<input>
<ID>IN_B_0</ID>374 </input>
<input>
<ID>IN_B_1</ID>380 </input>
<input>
<ID>IN_B_2</ID>402 </input>
<input>
<ID>IN_B_3</ID>408 </input>
<output>
<ID>OUT_0</ID>552 </output>
<output>
<ID>OUT_1</ID>551 </output>
<output>
<ID>OUT_2</ID>548 </output>
<output>
<ID>OUT_3</ID>522 </output>
<output>
<ID>carry_out</ID>553 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_FULLADDER_4BIT</type>
<position>84,-39</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>111 </input>
<input>
<ID>IN_2</ID>118 </input>
<input>
<ID>IN_3</ID>119 </input>
<input>
<ID>IN_B_0</ID>76 </input>
<input>
<ID>IN_B_1</ID>27 </input>
<input>
<ID>IN_B_2</ID>26 </input>
<input>
<ID>IN_B_3</ID>75 </input>
<output>
<ID>OUT_0</ID>59 </output>
<output>
<ID>OUT_1</ID>61 </output>
<output>
<ID>OUT_2</ID>60 </output>
<output>
<ID>OUT_3</ID>62 </output>
<output>
<ID>carry_out</ID>131 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>412</ID>
<type>AE_FULLADDER_4BIT</type>
<position>549.5,3.5</position>
<input>
<ID>IN_0</ID>424 </input>
<input>
<ID>IN_1</ID>423 </input>
<input>
<ID>IN_2</ID>422 </input>
<input>
<ID>IN_3</ID>417 </input>
<input>
<ID>IN_B_0</ID>410 </input>
<input>
<ID>IN_B_1</ID>411 </input>
<input>
<ID>IN_B_2</ID>412 </input>
<input>
<ID>IN_B_3</ID>414 </input>
<output>
<ID>OUT_0</ID>521 </output>
<output>
<ID>OUT_1</ID>519 </output>
<output>
<ID>OUT_2</ID>516 </output>
<output>
<ID>OUT_3</ID>481 </output>
<input>
<ID>carry_in</ID>553 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>413</ID>
<type>EE_VDD</type>
<position>533.5,-13.5</position>
<output>
<ID>OUT_0</ID>477 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_FULLADDER_4BIT</type>
<position>143,-26</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>210 </input>
<input>
<ID>IN_2</ID>209 </input>
<input>
<ID>IN_3</ID>216 </input>
<input>
<ID>IN_B_0</ID>59 </input>
<input>
<ID>IN_B_1</ID>61 </input>
<input>
<ID>IN_B_2</ID>60 </input>
<input>
<ID>IN_B_3</ID>62 </input>
<output>
<ID>OUT_0</ID>149 </output>
<output>
<ID>OUT_1</ID>148 </output>
<output>
<ID>OUT_2</ID>147 </output>
<output>
<ID>OUT_3</ID>146 </output>
<input>
<ID>carry_in</ID>260 </input>
<output>
<ID>carry_out</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>37</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>117,-42.5</position>
<output>
<ID>A_less_B</ID>151 </output>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_B_0</ID>59 </input>
<input>
<ID>IN_B_1</ID>61 </input>
<input>
<ID>IN_B_2</ID>60 </input>
<input>
<ID>IN_B_3</ID>62 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>39</ID>
<type>EE_VDD</type>
<position>107,-47.5</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>EE_VDD</type>
<position>107.5,-44.5</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>41</ID>
<type>AE_FULLADDER_4BIT</type>
<position>76,-75.5</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_3</ID>260 </input>
<input>
<ID>IN_B_0</ID>274 </input>
<input>
<ID>IN_B_1</ID>278 </input>
<input>
<ID>IN_B_2</ID>280 </input>
<input>
<ID>IN_B_3</ID>281 </input>
<output>
<ID>OUT_0</ID>263 </output>
<output>
<ID>OUT_1</ID>264 </output>
<output>
<ID>OUT_2</ID>262 </output>
<output>
<ID>OUT_3</ID>266 </output>
<input>
<ID>carry_in</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>53,-6.5</position>
<gparam>LABEL_TEXT is minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>61,-7</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>74.5,-6</position>
<gparam>LABEL_TEXT pressd minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AI_XOR2</type>
<position>-101.5,-25.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>421 </input>
<output>
<ID>OUT</ID>431 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AI_XOR2</type>
<position>62,-12</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>260 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AI_XOR2</type>
<position>-101.5,-29.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>420 </input>
<output>
<ID>OUT</ID>432 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_FULLADDER_4BIT</type>
<position>143,-63</position>
<input>
<ID>IN_0</ID>267 </input>
<input>
<ID>IN_1</ID>268 </input>
<input>
<ID>IN_2</ID>269 </input>
<input>
<ID>IN_3</ID>265 </input>
<input>
<ID>IN_B_0</ID>112 </input>
<input>
<ID>IN_B_1</ID>114 </input>
<input>
<ID>IN_B_2</ID>113 </input>
<input>
<ID>IN_B_3</ID>115 </input>
<output>
<ID>OUT_0</ID>157 </output>
<output>
<ID>OUT_1</ID>158 </output>
<output>
<ID>OUT_2</ID>159 </output>
<output>
<ID>OUT_3</ID>161 </output>
<input>
<ID>carry_in</ID>164 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>55</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>120.5,-78</position>
<output>
<ID>A_less_B</ID>162 </output>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_3</ID>116 </input>
<input>
<ID>IN_B_0</ID>112 </input>
<input>
<ID>IN_B_1</ID>114 </input>
<input>
<ID>IN_B_2</ID>113 </input>
<input>
<ID>IN_B_3</ID>115 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>61</ID>
<type>EE_VDD</type>
<position>115.5,-83</position>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>DD_KEYPAD_HEX</type>
<position>212,-38.5</position>
<output>
<ID>OUT_0</ID>35 </output>
<output>
<ID>OUT_1</ID>36 </output>
<output>
<ID>OUT_2</ID>37 </output>
<output>
<ID>OUT_3</ID>38 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>63</ID>
<type>GA_LED</type>
<position>166.5,-74.5</position>
<input>
<ID>N_in2</ID>121 </input>
<input>
<ID>N_in3</ID>207 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>DD_KEYPAD_HEX</type>
<position>185.5,-50.5</position>
<output>
<ID>OUT_0</ID>49 </output>
<output>
<ID>OUT_1</ID>48 </output>
<output>
<ID>OUT_2</ID>47 </output>
<output>
<ID>OUT_3</ID>46 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_FULLADDER_4BIT</type>
<position>240,-44</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>48 </input>
<input>
<ID>IN_2</ID>47 </input>
<input>
<ID>IN_3</ID>46 </input>
<input>
<ID>IN_B_0</ID>35 </input>
<input>
<ID>IN_B_1</ID>36 </input>
<input>
<ID>IN_B_2</ID>37 </input>
<input>
<ID>IN_B_3</ID>38 </input>
<output>
<ID>OUT_0</ID>39 </output>
<output>
<ID>OUT_1</ID>41 </output>
<output>
<ID>OUT_2</ID>40 </output>
<output>
<ID>OUT_3</ID>42 </output>
<output>
<ID>carry_out</ID>153 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>67</ID>
<type>AE_FULLADDER_4BIT</type>
<position>289,-31</position>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>50 </input>
<input>
<ID>IN_B_0</ID>39 </input>
<input>
<ID>IN_B_1</ID>41 </input>
<input>
<ID>IN_B_2</ID>40 </input>
<input>
<ID>IN_B_3</ID>42 </input>
<output>
<ID>OUT_0</ID>172 </output>
<output>
<ID>OUT_1</ID>171 </output>
<output>
<ID>OUT_2</ID>165 </output>
<output>
<ID>OUT_3</ID>156 </output>
<output>
<ID>carry_out</ID>201 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>70</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>165,-26.5</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>148 </input>
<input>
<ID>IN_2</ID>147 </input>
<input>
<ID>IN_3</ID>146 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_OR2</type>
<position>122.5,-47.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>208 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>166.5,-63.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>158 </input>
<input>
<ID>IN_2</ID>159 </input>
<input>
<ID>IN_3</ID>161 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_OR2</type>
<position>126,-89.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>296 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>277,-47.5</position>
<output>
<ID>A_less_B</ID>173 </output>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_3</ID>43 </input>
<input>
<ID>IN_B_0</ID>39 </input>
<input>
<ID>IN_B_1</ID>41 </input>
<input>
<ID>IN_B_2</ID>40 </input>
<input>
<ID>IN_B_3</ID>42 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>76</ID>
<type>EE_VDD</type>
<position>267,-52.5</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>77</ID>
<type>EE_VDD</type>
<position>267.5,-49.5</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>78</ID>
<type>AI_XOR2</type>
<position>112,-80</position>
<input>
<ID>IN_0</ID>166 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AI_XOR2</type>
<position>-101.5,-33.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>419 </input>
<output>
<ID>OUT</ID>433 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>EE_VDD</type>
<position>108,-79</position>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>166.5,-76.5</position>
<input>
<ID>N_in2</ID>123 </input>
<input>
<ID>N_in3</ID>121 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AI_XOR2</type>
<position>-101.5,-37.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>418 </input>
<output>
<ID>OUT</ID>434 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>DD_KEYPAD_HEX</type>
<position>212.5,-75</position>
<output>
<ID>OUT_0</ID>51 </output>
<output>
<ID>OUT_1</ID>53 </output>
<output>
<ID>OUT_2</ID>57 </output>
<output>
<ID>OUT_3</ID>58 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>DD_KEYPAD_HEX</type>
<position>188,-87</position>
<output>
<ID>OUT_0</ID>137 </output>
<output>
<ID>OUT_1</ID>127 </output>
<output>
<ID>OUT_2</ID>126 </output>
<output>
<ID>OUT_3</ID>125 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>85</ID>
<type>AE_FULLADDER_4BIT</type>
<position>240,-79.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>127 </input>
<input>
<ID>IN_2</ID>126 </input>
<input>
<ID>IN_3</ID>125 </input>
<input>
<ID>IN_B_0</ID>51 </input>
<input>
<ID>IN_B_1</ID>53 </input>
<input>
<ID>IN_B_2</ID>57 </input>
<input>
<ID>IN_B_3</ID>58 </input>
<output>
<ID>OUT_0</ID>74 </output>
<output>
<ID>OUT_1</ID>101 </output>
<output>
<ID>OUT_2</ID>98 </output>
<output>
<ID>OUT_3</ID>102 </output>
<input>
<ID>carry_in</ID>153 </input>
<output>
<ID>carry_out</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>86</ID>
<type>AE_FULLADDER_4BIT</type>
<position>291.5,-68</position>
<input>
<ID>IN_1</ID>150 </input>
<input>
<ID>IN_2</ID>150 </input>
<input>
<ID>IN_B_0</ID>74 </input>
<input>
<ID>IN_B_1</ID>101 </input>
<input>
<ID>IN_B_2</ID>98 </input>
<input>
<ID>IN_B_3</ID>102 </input>
<output>
<ID>OUT_0</ID>180 </output>
<output>
<ID>OUT_1</ID>182 </output>
<output>
<ID>OUT_2</ID>183 </output>
<output>
<ID>OUT_3</ID>184 </output>
<input>
<ID>carry_in</ID>201 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>92</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>280.5,-83</position>
<output>
<ID>A_less_B</ID>185 </output>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_3</ID>103 </input>
<input>
<ID>IN_B_0</ID>74 </input>
<input>
<ID>IN_B_1</ID>101 </input>
<input>
<ID>IN_B_2</ID>98 </input>
<input>
<ID>IN_B_3</ID>102 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>93</ID>
<type>EE_VDD</type>
<position>275.5,-88</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>114</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>302,-31</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>171 </input>
<input>
<ID>IN_2</ID>165 </input>
<input>
<ID>IN_3</ID>156 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 8</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_OR2</type>
<position>283.5,-53</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>303.5,-68.5</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>182 </input>
<input>
<ID>IN_2</ID>183 </input>
<input>
<ID>IN_3</ID>184 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_OR2</type>
<position>286,-94.5</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>200 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>AI_XOR2</type>
<position>272,-85</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>201 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>EE_VDD</type>
<position>268,-84</position>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>129</ID>
<type>GA_LED</type>
<position>166.5,-78.5</position>
<input>
<ID>N_in0</ID>163 </input>
<input>
<ID>N_in2</ID>163 </input>
<input>
<ID>N_in3</ID>123 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>FF_GND</type>
<position>-37,-29.5</position>
<output>
<ID>OUT_0</ID>403 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>173</ID>
<type>FF_GND</type>
<position>-37,-41.5</position>
<output>
<ID>OUT_0</ID>404 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>174</ID>
<type>GA_LED</type>
<position>166.5,-80.5</position>
<input>
<ID>N_in3</ID>163 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>FF_GND</type>
<position>-36.5,-65.5</position>
<output>
<ID>OUT_0</ID>406 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_AND2</type>
<position>82,-9.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>AI_XOR2</type>
<position>134.5,-27</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>219 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>190</ID>
<type>AI_XOR2</type>
<position>134.5,-31</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>AI_XOR2</type>
<position>134.5,-35</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>AI_XOR2</type>
<position>134.5,-39</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>221 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>193</ID>
<type>FF_GND</type>
<position>-36.5,-77.5</position>
<output>
<ID>OUT_0</ID>407 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>195</ID>
<type>AI_XOR2</type>
<position>66,-24</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>273 </input>
<output>
<ID>OUT</ID>259 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>198</ID>
<type>AI_XOR2</type>
<position>66,-28</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AI_XOR2</type>
<position>66,-32</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>271 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>AI_XOR2</type>
<position>66,-36</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>270 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>FF_GND</type>
<position>130.5,-28</position>
<output>
<ID>OUT_0</ID>219 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>202</ID>
<type>FF_GND</type>
<position>130.5,-40</position>
<output>
<ID>OUT_0</ID>221 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>203</ID>
<type>FF_GND</type>
<position>131,-64</position>
<output>
<ID>OUT_0</ID>252 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>204</ID>
<type>FF_GND</type>
<position>131,-76</position>
<output>
<ID>OUT_0</ID>253 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>206</ID>
<type>AI_XOR2</type>
<position>65,-65</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>291 </input>
<output>
<ID>OUT</ID>274 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>AI_XOR2</type>
<position>65,-69</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>290 </input>
<output>
<ID>OUT</ID>278 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>208</ID>
<type>AI_XOR2</type>
<position>65,-73</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>289 </input>
<output>
<ID>OUT</ID>280 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>209</ID>
<type>AI_XOR2</type>
<position>65,-77</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>288 </input>
<output>
<ID>OUT</ID>281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>AI_XOR2</type>
<position>135,-63</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>AI_XOR2</type>
<position>135,-67</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>AI_XOR2</type>
<position>135,-71</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>269 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>AI_XOR2</type>
<position>135,-75</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>253 </input>
<output>
<ID>OUT</ID>265 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>DD_KEYPAD_HEX</type>
<position>50.5,-74.5</position>
<output>
<ID>OUT_0</ID>291 </output>
<output>
<ID>OUT_1</ID>290 </output>
<output>
<ID>OUT_2</ID>289 </output>
<output>
<ID>OUT_3</ID>288 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>215</ID>
<type>AI_XOR2</type>
<position>-102.5,-66.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>429 </input>
<output>
<ID>OUT</ID>435 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>DD_KEYPAD_HEX</type>
<position>26,-88</position>
<output>
<ID>OUT_0</ID>105 </output>
<output>
<ID>OUT_1</ID>104 </output>
<output>
<ID>OUT_2</ID>96 </output>
<output>
<ID>OUT_3</ID>95 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>217</ID>
<type>AE_FULLADDER_4BIT</type>
<position>84,-79</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>104 </input>
<input>
<ID>IN_2</ID>96 </input>
<input>
<ID>IN_3</ID>95 </input>
<input>
<ID>IN_B_0</ID>263 </input>
<input>
<ID>IN_B_1</ID>264 </input>
<input>
<ID>IN_B_2</ID>262 </input>
<input>
<ID>IN_B_3</ID>266 </input>
<output>
<ID>OUT_0</ID>112 </output>
<output>
<ID>OUT_1</ID>114 </output>
<output>
<ID>OUT_2</ID>113 </output>
<output>
<ID>OUT_3</ID>115 </output>
<input>
<ID>carry_in</ID>131 </input>
<output>
<ID>carry_out</ID>296 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>218</ID>
<type>AI_XOR2</type>
<position>381.5,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>325 </input>
<output>
<ID>OUT</ID>279 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>AI_XOR2</type>
<position>385.5,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>326 </input>
<output>
<ID>OUT</ID>277 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>AI_XOR2</type>
<position>389.5,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>327 </input>
<output>
<ID>OUT</ID>276 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>AI_XOR2</type>
<position>393.5,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>328 </input>
<output>
<ID>OUT</ID>275 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>30,-28</position>
<gparam>LABEL_TEXT /</gparam>
<gparam>TEXT_HEIGHT 12</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>DD_KEYPAD_HEX</type>
<position>490,21.5</position>
<output>
<ID>OUT_0</ID>558 </output>
<output>
<ID>OUT_1</ID>557 </output>
<output>
<ID>OUT_2</ID>556 </output>
<output>
<ID>OUT_3</ID>555 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>224</ID>
<type>AI_XOR2</type>
<position>-102.5,-70.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>428 </input>
<output>
<ID>OUT</ID>436 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>AI_XOR2</type>
<position>-102.5,-74.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>427 </input>
<output>
<ID>OUT</ID>437 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>226</ID>
<type>AI_XOR2</type>
<position>-102.5,-78.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>426 </input>
<output>
<ID>OUT</ID>438 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>DD_KEYPAD_HEX</type>
<position>-115.5,-35</position>
<output>
<ID>OUT_0</ID>421 </output>
<output>
<ID>OUT_1</ID>420 </output>
<output>
<ID>OUT_2</ID>419 </output>
<output>
<ID>OUT_3</ID>418 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 4</lparam></gate>
<gate>
<ID>228</ID>
<type>AE_FULLADDER_4BIT</type>
<position>379.5,-15.5</position>
<input>
<ID>IN_1</ID>292 </input>
<input>
<ID>IN_3</ID>292 </input>
<input>
<ID>IN_B_0</ID>275 </input>
<input>
<ID>IN_B_1</ID>276 </input>
<input>
<ID>IN_B_2</ID>277 </input>
<input>
<ID>IN_B_3</ID>279 </input>
<output>
<ID>OUT_0</ID>297 </output>
<output>
<ID>OUT_1</ID>299 </output>
<output>
<ID>OUT_2</ID>295 </output>
<output>
<ID>OUT_3</ID>298 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>229</ID>
<type>AI_XOR2</type>
<position>-32.5,-64.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>406 </input>
<output>
<ID>OUT</ID>415 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_TOGGLE</type>
<position>-104.5,-8.5</position>
<output>
<ID>OUT_0</ID>284 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>231</ID>
<type>AI_XOR2</type>
<position>-32.5,-68.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>405 </input>
<output>
<ID>OUT</ID>416 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>232</ID>
<type>DD_KEYPAD_HEX</type>
<position>-142.5,-48.5</position>
<output>
<ID>OUT_0</ID>341 </output>
<output>
<ID>OUT_1</ID>344 </output>
<output>
<ID>OUT_2</ID>376 </output>
<output>
<ID>OUT_3</ID>377 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>233</ID>
<type>AI_XOR2</type>
<position>-32.5,-72.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>405 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>234</ID>
<type>AI_XOR2</type>
<position>-32.5,-76.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>407 </input>
<output>
<ID>OUT</ID>413 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>235</ID>
<type>DD_KEYPAD_HEX</type>
<position>-117,-76</position>
<output>
<ID>OUT_0</ID>429 </output>
<output>
<ID>OUT_1</ID>428 </output>
<output>
<ID>OUT_2</ID>427 </output>
<output>
<ID>OUT_3</ID>426 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>236</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-83.5,-40.5</position>
<input>
<ID>IN_0</ID>341 </input>
<input>
<ID>IN_1</ID>344 </input>
<input>
<ID>IN_2</ID>376 </input>
<input>
<ID>IN_3</ID>377 </input>
<input>
<ID>IN_B_0</ID>431 </input>
<input>
<ID>IN_B_1</ID>432 </input>
<input>
<ID>IN_B_2</ID>433 </input>
<input>
<ID>IN_B_3</ID>434 </input>
<output>
<ID>OUT_0</ID>287 </output>
<output>
<ID>OUT_1</ID>294 </output>
<output>
<ID>OUT_2</ID>293 </output>
<output>
<ID>OUT_3</ID>300 </output>
<input>
<ID>carry_in</ID>409 </input>
<output>
<ID>carry_out</ID>381 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>238</ID>
<type>DD_KEYPAD_HEX</type>
<position>-141.5,-89.5</position>
<output>
<ID>OUT_0</ID>320 </output>
<output>
<ID>OUT_1</ID>319 </output>
<output>
<ID>OUT_2</ID>309 </output>
<output>
<ID>OUT_3</ID>308 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>240</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-83.5,-80.5</position>
<input>
<ID>IN_0</ID>320 </input>
<input>
<ID>IN_1</ID>319 </input>
<input>
<ID>IN_2</ID>309 </input>
<input>
<ID>IN_3</ID>308 </input>
<input>
<ID>IN_B_0</ID>435 </input>
<input>
<ID>IN_B_1</ID>436 </input>
<input>
<ID>IN_B_2</ID>437 </input>
<input>
<ID>IN_B_3</ID>438 </input>
<output>
<ID>OUT_0</ID>354 </output>
<output>
<ID>OUT_1</ID>356 </output>
<output>
<ID>OUT_2</ID>355 </output>
<output>
<ID>OUT_3</ID>363 </output>
<input>
<ID>carry_in</ID>381 </input>
<output>
<ID>carry_out</ID>430 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_FULLADDER_4BIT</type>
<position>370.5,-29</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>331 </input>
<input>
<ID>IN_2</ID>330 </input>
<input>
<ID>IN_3</ID>329 </input>
<input>
<ID>IN_B_0</ID>297 </input>
<input>
<ID>IN_B_1</ID>299 </input>
<input>
<ID>IN_B_2</ID>295 </input>
<input>
<ID>IN_B_3</ID>298 </input>
<output>
<ID>OUT_0</ID>339 </output>
<output>
<ID>OUT_1</ID>338 </output>
<output>
<ID>OUT_2</ID>337 </output>
<output>
<ID>OUT_3</ID>340 </output>
<output>
<ID>carry_out</ID>357 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>242</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-24.5,-27.5</position>
<input>
<ID>IN_0</ID>400 </input>
<input>
<ID>IN_1</ID>399 </input>
<input>
<ID>IN_2</ID>398 </input>
<input>
<ID>IN_3</ID>401 </input>
<input>
<ID>IN_B_0</ID>287 </input>
<input>
<ID>IN_B_1</ID>294 </input>
<input>
<ID>IN_B_2</ID>293 </input>
<input>
<ID>IN_B_3</ID>300 </input>
<output>
<ID>OUT_0</ID>385 </output>
<output>
<ID>OUT_1</ID>384 </output>
<output>
<ID>OUT_2</ID>383 </output>
<output>
<ID>OUT_3</ID>382 </output>
<input>
<ID>carry_in</ID>409 </input>
<output>
<ID>carry_out</ID>393 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>244</ID>
<type>DD_KEYPAD_HEX</type>
<position>344,24.5</position>
<output>
<ID>OUT_0</ID>336 </output>
<output>
<ID>OUT_1</ID>335 </output>
<output>
<ID>OUT_2</ID>334 </output>
<output>
<ID>OUT_3</ID>333 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>245</ID>
<type>DD_KEYPAD_HEX</type>
<position>355.5,24.5</position>
<output>
<ID>OUT_0</ID>332 </output>
<output>
<ID>OUT_1</ID>331 </output>
<output>
<ID>OUT_2</ID>330 </output>
<output>
<ID>OUT_3</ID>329 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>246</ID>
<type>DD_KEYPAD_HEX</type>
<position>376.5,24.5</position>
<output>
<ID>OUT_0</ID>324 </output>
<output>
<ID>OUT_1</ID>323 </output>
<output>
<ID>OUT_2</ID>322 </output>
<output>
<ID>OUT_3</ID>321 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>248</ID>
<type>DD_KEYPAD_HEX</type>
<position>391,24</position>
<output>
<ID>OUT_0</ID>328 </output>
<output>
<ID>OUT_1</ID>327 </output>
<output>
<ID>OUT_2</ID>326 </output>
<output>
<ID>OUT_3</ID>325 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_LABEL</type>
<position>-137.5,-29.5</position>
<gparam>LABEL_TEXT /</gparam>
<gparam>TEXT_HEIGHT 12</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>GA_LED</type>
<position>276,6.5</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>-50.5,-44</position>
<output>
<ID>A_less_B</ID>386 </output>
<input>
<ID>IN_0</ID>302 </input>
<input>
<ID>IN_3</ID>301 </input>
<input>
<ID>IN_B_0</ID>287 </input>
<input>
<ID>IN_B_1</ID>294 </input>
<input>
<ID>IN_B_2</ID>293 </input>
<input>
<ID>IN_B_3</ID>300 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_TOGGLE</type>
<position>305.5,14</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>254</ID>
<type>EE_VDD</type>
<position>-60.5,-49</position>
<output>
<ID>OUT_0</ID>301 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>257</ID>
<type>CC_PULSE</type>
<position>355,38.5</position>
<output>
<ID>OUT_0</ID>306 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>EE_VDD</type>
<position>-60,-46</position>
<output>
<ID>OUT_0</ID>302 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>259</ID>
<type>BE_JKFF_LOW</type>
<position>360,38.5</position>
<input>
<ID>J</ID>306 </input>
<input>
<ID>K</ID>306 </input>
<output>
<ID>Q</ID>305 </output>
<input>
<ID>clock</ID>306 </input>
<output>
<ID>nQ</ID>292 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>260</ID>
<type>DD_KEYPAD_HEX</type>
<position>489.5,5</position>
<output>
<ID>OUT_0</ID>562 </output>
<output>
<ID>OUT_1</ID>561 </output>
<output>
<ID>OUT_2</ID>560 </output>
<output>
<ID>OUT_3</ID>559 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>261</ID>
<type>GA_LED</type>
<position>366.5,24.5</position>
<input>
<ID>N_in1</ID>307 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>-114.5,-8</position>
<gparam>LABEL_TEXT is minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>264</ID>
<type>GA_LED</type>
<position>366.5,22.5</position>
<input>
<ID>N_in2</ID>305 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>265</ID>
<type>AA_TOGGLE</type>
<position>-106.5,-8.5</position>
<output>
<ID>OUT_0</ID>283 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>266</ID>
<type>GA_LED</type>
<position>366.5,26.5</position>
<input>
<ID>N_in1</ID>305 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>AA_LABEL</type>
<position>-93,-7.5</position>
<gparam>LABEL_TEXT pressd minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>268</ID>
<type>GA_LED</type>
<position>368.5,24.5</position>
<input>
<ID>N_in1</ID>307 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>271</ID>
<type>AI_XOR2</type>
<position>-105.5,-13.5</position>
<input>
<ID>IN_0</ID>284 </input>
<input>
<ID>IN_1</ID>283 </input>
<output>
<ID>OUT</ID>409 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>272</ID>
<type>GA_LED</type>
<position>364.5,24.5</position>
<input>
<ID>N_in1</ID>307 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>273</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-24.5,-64.5</position>
<input>
<ID>IN_0</ID>415 </input>
<input>
<ID>IN_1</ID>416 </input>
<input>
<ID>IN_3</ID>413 </input>
<input>
<ID>IN_B_0</ID>354 </input>
<input>
<ID>IN_B_1</ID>356 </input>
<input>
<ID>IN_B_2</ID>355 </input>
<input>
<ID>IN_B_3</ID>363 </input>
<output>
<ID>OUT_0</ID>387 </output>
<output>
<ID>OUT_1</ID>388 </output>
<output>
<ID>OUT_2</ID>389 </output>
<output>
<ID>OUT_3</ID>390 </output>
<input>
<ID>carry_in</ID>393 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>274</ID>
<type>AE_OR2</type>
<position>366.5,34.5</position>
<input>
<ID>IN_0</ID>305 </input>
<input>
<ID>IN_1</ID>292 </input>
<output>
<ID>OUT</ID>307 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>-47,-79.5</position>
<output>
<ID>A_less_B</ID>391 </output>
<input>
<ID>IN_0</ID>395 </input>
<input>
<ID>IN_3</ID>375 </input>
<input>
<ID>IN_B_0</ID>354 </input>
<input>
<ID>IN_B_1</ID>356 </input>
<input>
<ID>IN_B_2</ID>355 </input>
<input>
<ID>IN_B_3</ID>363 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_LABEL</type>
<position>409,4.5</position>
<gparam>LABEL_TEXT minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>277</ID>
<type>AI_XOR2</type>
<position>350,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>321 </input>
<output>
<ID>OUT</ID>313 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>AI_XOR2</type>
<position>354,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>312 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>AI_XOR2</type>
<position>358,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>323 </input>
<output>
<ID>OUT</ID>311 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>670</ID>
<type>BB_CLOCK</type>
<position>491.5,-23</position>
<output>
<ID>CLK</ID>303 </output>
<gparam>angle 0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>281</ID>
<type>AI_XOR2</type>
<position>362,-1</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>324 </input>
<output>
<ID>OUT</ID>310 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>AE_FULLADDER_4BIT</type>
<position>348,-15.5</position>
<input>
<ID>IN_1</ID>292 </input>
<input>
<ID>IN_3</ID>292 </input>
<input>
<ID>IN_B_0</ID>310 </input>
<input>
<ID>IN_B_1</ID>311 </input>
<input>
<ID>IN_B_2</ID>312 </input>
<input>
<ID>IN_B_3</ID>313 </input>
<output>
<ID>OUT_0</ID>316 </output>
<output>
<ID>OUT_1</ID>318 </output>
<output>
<ID>OUT_2</ID>315 </output>
<output>
<ID>OUT_3</ID>317 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>672</ID>
<type>CC_PULSE</type>
<position>518,-20</position>
<output>
<ID>OUT_0</ID>261 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>283</ID>
<type>AE_FULLADDER_4BIT</type>
<position>339,-29</position>
<input>
<ID>IN_0</ID>336 </input>
<input>
<ID>IN_1</ID>335 </input>
<input>
<ID>IN_2</ID>334 </input>
<input>
<ID>IN_3</ID>333 </input>
<input>
<ID>IN_B_0</ID>316 </input>
<input>
<ID>IN_B_1</ID>318 </input>
<input>
<ID>IN_B_2</ID>315 </input>
<input>
<ID>IN_B_3</ID>317 </input>
<output>
<ID>OUT_0</ID>347 </output>
<output>
<ID>OUT_1</ID>346 </output>
<output>
<ID>OUT_2</ID>345 </output>
<output>
<ID>OUT_3</ID>348 </output>
<input>
<ID>carry_in</ID>357 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>673</ID>
<type>CC_PULSE</type>
<position>515,-34.5</position>
<output>
<ID>OUT_0</ID>554 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>284</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>359.5,-44.5</position>
<output>
<ID>A_less_B</ID>549 </output>
<input>
<ID>IN_0</ID>343 </input>
<input>
<ID>IN_3</ID>342 </input>
<input>
<ID>IN_B_0</ID>339 </input>
<input>
<ID>IN_B_1</ID>338 </input>
<input>
<ID>IN_B_2</ID>337 </input>
<input>
<ID>IN_B_3</ID>340 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>285</ID>
<type>EE_VDD</type>
<position>-52,-84.5</position>
<output>
<ID>OUT_0</ID>375 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>286</ID>
<type>EE_VDD</type>
<position>354.5,-39.5</position>
<output>
<ID>OUT_0</ID>342 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>287</ID>
<type>EE_VDD</type>
<position>357.5,-39.5</position>
<output>
<ID>OUT_0</ID>343 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>288</ID>
<type>AE_FULLADDER_4BIT</type>
<position>367,-53</position>
<input>
<ID>IN_1</ID>358 </input>
<input>
<ID>IN_2</ID>358 </input>
<input>
<ID>IN_B_0</ID>339 </input>
<input>
<ID>IN_B_1</ID>338 </input>
<input>
<ID>IN_B_2</ID>337 </input>
<input>
<ID>IN_B_3</ID>340 </input>
<output>
<ID>OUT_0</ID>367 </output>
<output>
<ID>OUT_1</ID>366 </output>
<output>
<ID>OUT_2</ID>365 </output>
<output>
<ID>OUT_3</ID>364 </output>
<output>
<ID>carry_out</ID>550 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>290</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>328,-44</position>
<output>
<ID>A_less_B</ID>352 </output>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_3</ID>349 </input>
<input>
<ID>IN_B_0</ID>347 </input>
<input>
<ID>IN_B_1</ID>346 </input>
<input>
<ID>IN_B_2</ID>345 </input>
<input>
<ID>IN_B_3</ID>348 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>295</ID>
<type>EE_VDD</type>
<position>323,-39</position>
<output>
<ID>OUT_0</ID>349 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>297</ID>
<type>AE_FULLADDER_4BIT</type>
<position>335.5,-53</position>
<input>
<ID>IN_1</ID>352 </input>
<input>
<ID>IN_2</ID>352 </input>
<input>
<ID>IN_B_0</ID>347 </input>
<input>
<ID>IN_B_1</ID>346 </input>
<input>
<ID>IN_B_2</ID>345 </input>
<input>
<ID>IN_B_3</ID>348 </input>
<output>
<ID>OUT_0</ID>542 </output>
<output>
<ID>OUT_1</ID>543 </output>
<output>
<ID>OUT_2</ID>544 </output>
<output>
<ID>OUT_3</ID>545 </output>
<input>
<ID>carry_in</ID>550 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>298</ID>
<type>AI_XOR2</type>
<position>359.5,-63</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>362 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>299</ID>
<type>AI_XOR2</type>
<position>363.5,-63</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>365 </input>
<output>
<ID>OUT</ID>361 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>300</ID>
<type>AI_XOR2</type>
<position>367.5,-63</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>360 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>301</ID>
<type>AI_XOR2</type>
<position>371.5,-63</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>367 </input>
<output>
<ID>OUT</ID>359 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>AE_FULLADDER_4BIT</type>
<position>360.5,-74</position>
<input>
<ID>IN_1</ID>353 </input>
<input>
<ID>IN_3</ID>353 </input>
<input>
<ID>IN_B_0</ID>359 </input>
<input>
<ID>IN_B_1</ID>360 </input>
<input>
<ID>IN_B_2</ID>361 </input>
<input>
<ID>IN_B_3</ID>362 </input>
<output>
<ID>OUT_0</ID>529 </output>
<output>
<ID>OUT_1</ID>528 </output>
<output>
<ID>OUT_2</ID>527 </output>
<output>
<ID>OUT_3</ID>526 </output>
<input>
<ID>carry_in</ID>358 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>304</ID>
<type>GA_LED</type>
<position>-1,-76</position>
<input>
<ID>N_in2</ID>378 </input>
<input>
<ID>N_in3</ID>396 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>305</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-2.5,-28</position>
<input>
<ID>IN_0</ID>385 </input>
<input>
<ID>IN_1</ID>384 </input>
<input>
<ID>IN_2</ID>383 </input>
<input>
<ID>IN_3</ID>382 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_OR2</type>
<position>-45,-49</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>439 </input>
<output>
<ID>OUT</ID>397 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>AE_SMALL_INVERTER</type>
<position>349,-56.5</position>
<input>
<ID>IN_0</ID>358 </input>
<output>
<ID>OUT_0</ID>353 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>308</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>367,-83.5</position>
<input>
<ID>IN_0</ID>529 </input>
<input>
<ID>IN_1</ID>528 </input>
<input>
<ID>IN_2</ID>527 </input>
<input>
<ID>IN_3</ID>526 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>309</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-1,-65</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>388 </input>
<input>
<ID>IN_2</ID>389 </input>
<input>
<ID>IN_3</ID>390 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 12</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>310</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>589,-37.5</position>
<input>
<ID>IN_0</ID>552 </input>
<input>
<ID>IN_1</ID>551 </input>
<input>
<ID>IN_2</ID>548 </input>
<input>
<ID>IN_3</ID>522 </input>
<input>
<ID>IN_4</ID>521 </input>
<input>
<ID>IN_5</ID>519 </input>
<input>
<ID>IN_6</ID>516 </input>
<input>
<ID>IN_7</ID>481 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>311</ID>
<type>AE_REGISTER8</type>
<position>534,-22</position>
<input>
<ID>IN_0</ID>552 </input>
<input>
<ID>IN_1</ID>551 </input>
<input>
<ID>IN_2</ID>548 </input>
<input>
<ID>IN_3</ID>522 </input>
<input>
<ID>IN_4</ID>521 </input>
<input>
<ID>IN_5</ID>519 </input>
<input>
<ID>IN_6</ID>516 </input>
<input>
<ID>IN_7</ID>481 </input>
<output>
<ID>OUT_0</ID>442 </output>
<output>
<ID>OUT_1</ID>441 </output>
<output>
<ID>OUT_2</ID>440 </output>
<output>
<ID>OUT_3</ID>425 </output>
<output>
<ID>OUT_4</ID>424 </output>
<output>
<ID>OUT_5</ID>423 </output>
<output>
<ID>OUT_6</ID>422 </output>
<output>
<ID>OUT_7</ID>417 </output>
<input>
<ID>clear</ID>554 </input>
<input>
<ID>clock</ID>303 </input>
<input>
<ID>load</ID>477 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>312</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>511,27</position>
<input>
<ID>IN_0</ID>555 </input>
<input>
<ID>IN_1</ID>556 </input>
<input>
<ID>IN_2</ID>557 </input>
<input>
<ID>IN_3</ID>558 </input>
<output>
<ID>carry_out</ID>373 </output>
<input>
<ID>clear</ID>554 </input>
<input>
<ID>clock</ID>303 </input>
<input>
<ID>load</ID>261 </input>
<input>
<ID>shift_enable</ID>769 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>313</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>510,10</position>
<input>
<ID>IN_0</ID>562 </input>
<input>
<ID>IN_1</ID>561 </input>
<input>
<ID>IN_2</ID>560 </input>
<input>
<ID>IN_3</ID>559 </input>
<output>
<ID>OUT_0</ID>372 </output>
<output>
<ID>OUT_1</ID>371 </output>
<output>
<ID>OUT_2</ID>370 </output>
<output>
<ID>OUT_3</ID>369 </output>
<output>
<ID>carry_out</ID>304 </output>
<input>
<ID>clear</ID>554 </input>
<input>
<ID>clock</ID>303 </input>
<input>
<ID>load</ID>261 </input>
<input>
<ID>shift_enable</ID>768 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>314</ID>
<type>AE_OR2</type>
<position>-42,-91</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>430 </input>
<output>
<ID>OUT</ID>443 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>315</ID>
<type>AI_XOR2</type>
<position>-55.5,-81.5</position>
<input>
<ID>IN_0</ID>394 </input>
<input>
<ID>IN_1</ID>393 </input>
<output>
<ID>OUT</ID>395 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>316</ID>
<type>EE_VDD</type>
<position>-59.5,-80.5</position>
<output>
<ID>OUT_0</ID>394 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>317</ID>
<type>GA_LED</type>
<position>-1,-78</position>
<input>
<ID>N_in2</ID>379 </input>
<input>
<ID>N_in3</ID>378 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>318</ID>
<type>GA_LED</type>
<position>-1,-80</position>
<input>
<ID>N_in0</ID>392 </input>
<input>
<ID>N_in2</ID>392 </input>
<input>
<ID>N_in3</ID>379 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>319</ID>
<type>GA_LED</type>
<position>-1,-82</position>
<input>
<ID>N_in3</ID>392 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>320</ID>
<type>AA_AND2</type>
<position>-85.5,-11</position>
<input>
<ID>IN_0</ID>283 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>396 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>321</ID>
<type>AI_XOR2</type>
<position>-33,-28.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>403 </input>
<output>
<ID>OUT</ID>400 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>322</ID>
<type>AI_XOR2</type>
<position>-33,-32.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>399 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>323</ID>
<type>AI_XOR2</type>
<position>-33,-36.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>398 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>324</ID>
<type>AI_XOR2</type>
<position>-33,-40.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>404 </input>
<output>
<ID>OUT</ID>401 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>325</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>510,-6</position>
<output>
<ID>OUT_0</ID>368 </output>
<output>
<ID>OUT_1</ID>351 </output>
<output>
<ID>OUT_2</ID>350 </output>
<output>
<ID>OUT_3</ID>314 </output>
<input>
<ID>carry_in</ID>304 </input>
<input>
<ID>clear</ID>554 </input>
<input>
<ID>clock</ID>303 </input>
<input>
<ID>load</ID>261 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>326</ID>
<type>AI_XOR2</type>
<position>-72.5,-54</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>381 </input>
<output>
<ID>OUT</ID>439 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>AI_XOR2</type>
<position>-36,-84.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>443 </input>
<output>
<ID>OUT</ID>405 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>330</ID>
<type>FF_GND</type>
<position>-198,-79.5</position>
<output>
<ID>OUT_0</ID>492 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>331</ID>
<type>AI_XOR2</type>
<position>-264,-68.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>505 </input>
<output>
<ID>OUT</ID>511 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>332</ID>
<type>AI_XOR2</type>
<position>-264,-72.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>504 </input>
<output>
<ID>OUT</ID>512 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>333</ID>
<type>AI_XOR2</type>
<position>-264,-76.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>503 </input>
<output>
<ID>OUT</ID>513 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>334</ID>
<type>AI_XOR2</type>
<position>-264,-80.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>514 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>335</ID>
<type>DD_KEYPAD_HEX</type>
<position>-277,-37</position>
<output>
<ID>OUT_0</ID>501 </output>
<output>
<ID>OUT_1</ID>500 </output>
<output>
<ID>OUT_2</ID>499 </output>
<output>
<ID>OUT_3</ID>498 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>336</ID>
<type>AI_XOR2</type>
<position>-194,-66.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>491 </input>
<output>
<ID>OUT</ID>495 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>337</ID>
<type>AA_TOGGLE</type>
<position>-266,-10.5</position>
<output>
<ID>OUT_0</ID>445 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>338</ID>
<type>AI_XOR2</type>
<position>-194,-70.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>490 </input>
<output>
<ID>OUT</ID>496 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>339</ID>
<type>DD_KEYPAD_HEX</type>
<position>-303.5,-54</position>
<output>
<ID>OUT_0</ID>456 </output>
<output>
<ID>OUT_1</ID>457 </output>
<output>
<ID>OUT_2</ID>463 </output>
<output>
<ID>OUT_3</ID>464 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>340</ID>
<type>AI_XOR2</type>
<position>-194,-74.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>490 </input>
<output>
<ID>OUT</ID>497 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>AI_XOR2</type>
<position>-194,-78.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>494 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>342</ID>
<type>DD_KEYPAD_HEX</type>
<position>-278.5,-78</position>
<output>
<ID>OUT_0</ID>505 </output>
<output>
<ID>OUT_1</ID>504 </output>
<output>
<ID>OUT_2</ID>503 </output>
<output>
<ID>OUT_3</ID>502 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>343</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-245,-42.5</position>
<input>
<ID>IN_0</ID>456 </input>
<input>
<ID>IN_1</ID>457 </input>
<input>
<ID>IN_2</ID>463 </input>
<input>
<ID>IN_3</ID>464 </input>
<input>
<ID>IN_B_0</ID>507 </input>
<input>
<ID>IN_B_1</ID>508 </input>
<input>
<ID>IN_B_2</ID>509 </input>
<input>
<ID>IN_B_3</ID>510 </input>
<output>
<ID>OUT_0</ID>446 </output>
<output>
<ID>OUT_1</ID>448 </output>
<output>
<ID>OUT_2</ID>447 </output>
<output>
<ID>OUT_3</ID>449 </output>
<input>
<ID>carry_in</ID>493 </input>
<output>
<ID>carry_out</ID>467 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>344</ID>
<type>DD_KEYPAD_HEX</type>
<position>-303,-91.5</position>
<output>
<ID>OUT_0</ID>455 </output>
<output>
<ID>OUT_1</ID>454 </output>
<output>
<ID>OUT_2</ID>453 </output>
<output>
<ID>OUT_3</ID>452 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>345</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-245,-82.5</position>
<input>
<ID>IN_0</ID>455 </input>
<input>
<ID>IN_1</ID>454 </input>
<input>
<ID>IN_2</ID>453 </input>
<input>
<ID>IN_3</ID>452 </input>
<input>
<ID>IN_B_0</ID>511 </input>
<input>
<ID>IN_B_1</ID>512 </input>
<input>
<ID>IN_B_2</ID>513 </input>
<input>
<ID>IN_B_3</ID>514 </input>
<output>
<ID>OUT_0</ID>458 </output>
<output>
<ID>OUT_1</ID>460 </output>
<output>
<ID>OUT_2</ID>459 </output>
<output>
<ID>OUT_3</ID>461 </output>
<input>
<ID>carry_in</ID>525 </input>
<output>
<ID>carry_out</ID>506 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>346</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-186,-29.5</position>
<input>
<ID>IN_0</ID>486 </input>
<input>
<ID>IN_1</ID>485 </input>
<input>
<ID>IN_2</ID>484 </input>
<input>
<ID>IN_3</ID>487 </input>
<input>
<ID>IN_B_0</ID>446 </input>
<input>
<ID>IN_B_1</ID>448 </input>
<input>
<ID>IN_B_2</ID>447 </input>
<input>
<ID>IN_B_3</ID>449 </input>
<output>
<ID>OUT_0</ID>471 </output>
<output>
<ID>OUT_1</ID>470 </output>
<output>
<ID>OUT_2</ID>469 </output>
<output>
<ID>OUT_3</ID>468 </output>
<input>
<ID>carry_in</ID>493 </input>
<output>
<ID>carry_out</ID>479 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>347</ID>
<type>AI_XOR2</type>
<position>-263,-27.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>348</ID>
<type>AI_XOR2</type>
<position>-263,-31.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>500 </input>
<output>
<ID>OUT</ID>508 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>349</ID>
<type>AA_LABEL</type>
<position>-299,-31.5</position>
<gparam>LABEL_TEXT /</gparam>
<gparam>TEXT_HEIGHT 12</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>-212,-46</position>
<output>
<ID>A_less_B</ID>472 </output>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_3</ID>450 </input>
<input>
<ID>IN_B_0</ID>446 </input>
<input>
<ID>IN_B_1</ID>448 </input>
<input>
<ID>IN_B_2</ID>447 </input>
<input>
<ID>IN_B_3</ID>449 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>351</ID>
<type>EE_VDD</type>
<position>-222,-51</position>
<output>
<ID>OUT_0</ID>450 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>352</ID>
<type>EE_VDD</type>
<position>-221.5,-48</position>
<output>
<ID>OUT_0</ID>451 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>353</ID>
<type>AA_LABEL</type>
<position>-276,-10</position>
<gparam>LABEL_TEXT is minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>354</ID>
<type>AA_TOGGLE</type>
<position>-268,-10.5</position>
<output>
<ID>OUT_0</ID>444 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_LABEL</type>
<position>-254.5,-9.5</position>
<gparam>LABEL_TEXT pressd minus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>356</ID>
<type>AI_XOR2</type>
<position>-267,-15.5</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>444 </input>
<output>
<ID>OUT</ID>493 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>AI_XOR2</type>
<position>-263,-35.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>499 </input>
<output>
<ID>OUT</ID>509 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>358</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-186,-66.5</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>496 </input>
<input>
<ID>IN_2</ID>497 </input>
<input>
<ID>IN_3</ID>494 </input>
<input>
<ID>IN_B_0</ID>458 </input>
<input>
<ID>IN_B_1</ID>460 </input>
<input>
<ID>IN_B_2</ID>459 </input>
<input>
<ID>IN_B_3</ID>461 </input>
<output>
<ID>OUT_0</ID>473 </output>
<output>
<ID>OUT_1</ID>474 </output>
<output>
<ID>OUT_2</ID>475 </output>
<output>
<ID>OUT_3</ID>476 </output>
<input>
<ID>carry_in</ID>479 </input>
<output>
<ID>carry_out</ID>520 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>359</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>-210,-81.5</position>
<output>
<ID>A_less_B</ID>523 </output>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_3</ID>462 </input>
<input>
<ID>IN_B_0</ID>458 </input>
<input>
<ID>IN_B_1</ID>460 </input>
<input>
<ID>IN_B_2</ID>459 </input>
<input>
<ID>IN_B_3</ID>461 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>360</ID>
<type>AI_XOR2</type>
<position>-263,-39.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>498 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>EE_VDD</type>
<position>-215.5,-86.5</position>
<output>
<ID>OUT_0</ID>462 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>362</ID>
<type>GA_LED</type>
<position>-162.5,-78</position>
<input>
<ID>N_in2</ID>465 </input>
<input>
<ID>N_in3</ID>482 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>363</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-164,-30</position>
<input>
<ID>IN_0</ID>471 </input>
<input>
<ID>IN_1</ID>470 </input>
<input>
<ID>IN_2</ID>469 </input>
<input>
<ID>IN_3</ID>468 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>364</ID>
<type>AE_OR2</type>
<position>-206.5,-51</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>515 </input>
<output>
<ID>OUT</ID>483 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>365</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-162.5,-67</position>
<input>
<ID>IN_0</ID>473 </input>
<input>
<ID>IN_1</ID>474 </input>
<input>
<ID>IN_2</ID>475 </input>
<input>
<ID>IN_3</ID>476 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>366</ID>
<type>AE_OR2</type>
<position>-203.5,-97.5</position>
<input>
<ID>IN_0</ID>523 </input>
<input>
<ID>IN_1</ID>506 </input>
<output>
<ID>OUT</ID>518 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>367</ID>
<type>AI_XOR2</type>
<position>-217,-83.5</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>479 </input>
<output>
<ID>OUT</ID>517 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>368</ID>
<type>EE_VDD</type>
<position>-221,-82.5</position>
<output>
<ID>OUT_0</ID>480 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>369</ID>
<type>GA_LED</type>
<position>-162.5,-80</position>
<input>
<ID>N_in0</ID>524 </input>
<input>
<ID>N_in2</ID>466 </input>
<input>
<ID>N_in3</ID>465 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>370</ID>
<type>GA_LED</type>
<position>-162.5,-82</position>
<input>
<ID>N_in0</ID>478 </input>
<input>
<ID>N_in2</ID>478 </input>
<input>
<ID>N_in3</ID>466 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>371</ID>
<type>GA_LED</type>
<position>-162.5,-84</position>
<input>
<ID>N_in1</ID>524 </input>
<input>
<ID>N_in3</ID>478 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>372</ID>
<type>AA_AND2</type>
<position>-247,-13</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>445 </input>
<output>
<ID>OUT</ID>482 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>373</ID>
<type>AI_XOR2</type>
<position>-194.5,-30.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>488 </input>
<output>
<ID>OUT</ID>486 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>AI_XOR2</type>
<position>-194.5,-34.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>483 </input>
<output>
<ID>OUT</ID>485 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>AI_XOR2</type>
<position>-194.5,-38.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>483 </input>
<output>
<ID>OUT</ID>484 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>376</ID>
<type>AI_XOR2</type>
<position>-194.5,-42.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>489 </input>
<output>
<ID>OUT</ID>487 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>377</ID>
<type>AI_XOR2</type>
<position>-234,-56</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>467 </input>
<output>
<ID>OUT</ID>515 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>378</ID>
<type>AI_XOR2</type>
<position>-199.5,-92.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>518 </input>
<output>
<ID>OUT</ID>490 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>FF_GND</type>
<position>-198.5,-31.5</position>
<output>
<ID>OUT_0</ID>488 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>380</ID>
<type>FF_GND</type>
<position>-198.5,-43.5</position>
<output>
<ID>OUT_0</ID>489 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>381</ID>
<type>FF_GND</type>
<position>-198,-67.5</position>
<output>
<ID>OUT_0</ID>491 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>382</ID>
<type>AE_SMALL_INVERTER</type>
<position>510,1</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>383</ID>
<type>AE_SMALL_INVERTER</type>
<position>509.5,18</position>
<input>
<ID>IN_0</ID>261 </input>
<output>
<ID>OUT_0</ID>768 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>384</ID>
<type>AE_SMALL_INVERTER</type>
<position>510,35</position>
<input>
<ID>IN_0</ID>261 </input>
<output>
<ID>OUT_0</ID>769 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>385</ID>
<type>GA_LED</type>
<position>-172,-78.5</position>
<input>
<ID>N_in3</ID>520 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>386</ID>
<type>AE_OR2</type>
<position>-245,-70</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>467 </input>
<output>
<ID>OUT</ID>525 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>387</ID>
<type>AI_XOR2</type>
<position>326,-63</position>
<input>
<ID>IN_0</ID>530 </input>
<input>
<ID>IN_1</ID>545 </input>
<output>
<ID>OUT</ID>534 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>388</ID>
<type>AI_XOR2</type>
<position>330,-63</position>
<input>
<ID>IN_0</ID>530 </input>
<input>
<ID>IN_1</ID>544 </input>
<output>
<ID>OUT</ID>533 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>769</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,32.5,510,33</points>
<connection>
<GID>384</GID>
<name>OUT_0</name></connection>
<intersection>32.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>511,32,511,32.5</points>
<connection>
<GID>312</GID>
<name>shift_enable</name></connection>
<intersection>32.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>510,32.5,511,32.5</points>
<intersection>510 0</intersection>
<intersection>511 1</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-9,61,-8.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-8.5,79,-8.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-10.5,63,-9</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-10.5,79,-10.5</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-36,80,-36</points>
<connection>
<GID>14</GID>
<name>OUT_2</name></connection>
<connection>
<GID>22</GID>
<name>IN_B_2</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-35,80,-35</points>
<connection>
<GID>14</GID>
<name>OUT_1</name></connection>
<connection>
<GID>22</GID>
<name>IN_B_1</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-41.5,226.5,-39</points>
<intersection>-41.5 3</intersection>
<intersection>-39 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-41.5,226.5,-41.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-39,236,-39</points>
<connection>
<GID>66</GID>
<name>IN_B_0</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-40,226.5,-39.5</points>
<intersection>-40 6</intersection>
<intersection>-39.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>217,-39.5,226.5,-39.5</points>
<connection>
<GID>62</GID>
<name>OUT_1</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>226.5,-40,236,-40</points>
<connection>
<GID>66</GID>
<name>IN_B_1</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-41,226.5,-37.5</points>
<intersection>-41 4</intersection>
<intersection>-37.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-37.5,226.5,-37.5</points>
<connection>
<GID>62</GID>
<name>OUT_2</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-41,236,-41</points>
<connection>
<GID>66</GID>
<name>IN_B_2</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-42,226.5,-35.5</points>
<intersection>-42 4</intersection>
<intersection>-35.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-35.5,226.5,-35.5</points>
<connection>
<GID>62</GID>
<name>OUT_3</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-42,236,-42</points>
<connection>
<GID>66</GID>
<name>IN_B_3</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-42.5,273,-42.5</points>
<connection>
<GID>75</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>252.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>252.5,-42.5,252.5,-26</points>
<intersection>-42.5 1</intersection>
<intersection>-26 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>252.5,-26,285,-26</points>
<connection>
<GID>67</GID>
<name>IN_B_0</name></connection>
<intersection>252.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-44.5,273,-44.5</points>
<connection>
<GID>75</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>66</GID>
<name>OUT_2</name></connection>
<intersection>254.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>254.5,-44.5,254.5,-28</points>
<intersection>-44.5 1</intersection>
<intersection>-28 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>254.5,-28,285,-28</points>
<connection>
<GID>67</GID>
<name>IN_B_2</name></connection>
<intersection>254.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-43.5,273,-43.5</points>
<connection>
<GID>75</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>66</GID>
<name>OUT_1</name></connection>
<intersection>253.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>253.5,-43.5,253.5,-27</points>
<intersection>-43.5 1</intersection>
<intersection>-27 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>253.5,-27,285,-27</points>
<connection>
<GID>67</GID>
<name>IN_B_1</name></connection>
<intersection>253.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-45.5,273,-45.5</points>
<connection>
<GID>75</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>66</GID>
<name>OUT_3</name></connection>
<intersection>256 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>256,-45.5,256,-29</points>
<intersection>-45.5 1</intersection>
<intersection>-29 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>256,-29,285,-29</points>
<connection>
<GID>67</GID>
<name>IN_B_3</name></connection>
<intersection>256 6</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>268,-52.5,273,-52.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<connection>
<GID>75</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>268.5,-49.5,273,-49.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<connection>
<GID>75</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-49,213,-47.5</points>
<intersection>-49 4</intersection>
<intersection>-47.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>190.5,-47.5,213,-47.5</points>
<connection>
<GID>64</GID>
<name>OUT_3</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>213,-49,236,-49</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-49.5,213,-48</points>
<intersection>-49.5 3</intersection>
<intersection>-48 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>190.5,-49.5,213,-49.5</points>
<connection>
<GID>64</GID>
<name>OUT_2</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>213,-48,236,-48</points>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-51.5,213,-47</points>
<intersection>-51.5 3</intersection>
<intersection>-47 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>190.5,-51.5,213,-51.5</points>
<connection>
<GID>64</GID>
<name>OUT_1</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>213,-47,236,-47</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-53.5,213,-46</points>
<intersection>-53.5 3</intersection>
<intersection>-46 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>190.5,-53.5,213,-53.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>213,-46,236,-46</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>283.5,-50,283.5,-34</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>-35 30</intersection>
<intersection>-34 31</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>283.5,-35,285,-35</points>
<connection>
<GID>67</GID>
<name>IN_2</name></connection>
<intersection>283.5 2</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>283.5,-34,285,-34</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>283.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-78,226.5,-74.5</points>
<intersection>-78 3</intersection>
<intersection>-74.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217.5,-78,226.5,-78</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-74.5,236,-74.5</points>
<connection>
<GID>85</GID>
<name>IN_B_0</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-76,226.5,-75.5</points>
<intersection>-76 7</intersection>
<intersection>-75.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>217.5,-76,226.5,-76</points>
<connection>
<GID>83</GID>
<name>OUT_1</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>226.5,-75.5,236,-75.5</points>
<connection>
<GID>85</GID>
<name>IN_B_1</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-76.5,226.5,-74</points>
<intersection>-76.5 4</intersection>
<intersection>-74 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217.5,-74,226.5,-74</points>
<connection>
<GID>83</GID>
<name>OUT_2</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-76.5,236,-76.5</points>
<connection>
<GID>85</GID>
<name>IN_B_2</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-77.5,226.5,-72</points>
<intersection>-77.5 4</intersection>
<intersection>-72 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217.5,-72,226.5,-72</points>
<connection>
<GID>83</GID>
<name>OUT_3</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-77.5,236,-77.5</points>
<connection>
<GID>85</GID>
<name>IN_B_3</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-37.5,113,-37.5</points>
<connection>
<GID>37</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>92.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>92.5,-37.5,92.5,-21</points>
<intersection>-37.5 1</intersection>
<intersection>-21 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>92.5,-21,139,-21</points>
<connection>
<GID>27</GID>
<name>IN_B_0</name></connection>
<intersection>92.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-39.5,113,-39.5</points>
<connection>
<GID>37</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>22</GID>
<name>OUT_2</name></connection>
<intersection>94.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>94.5,-39.5,94.5,-23</points>
<intersection>-39.5 1</intersection>
<intersection>-23 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>94.5,-23,139,-23</points>
<connection>
<GID>27</GID>
<name>IN_B_2</name></connection>
<intersection>94.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-38.5,113,-38.5</points>
<connection>
<GID>37</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>22</GID>
<name>OUT_1</name></connection>
<intersection>93.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>93.5,-38.5,93.5,-22</points>
<intersection>-38.5 1</intersection>
<intersection>-22 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>93.5,-22,139,-22</points>
<connection>
<GID>27</GID>
<name>IN_B_1</name></connection>
<intersection>93.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-40.5,113,-40.5</points>
<connection>
<GID>37</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>22</GID>
<name>OUT_3</name></connection>
<intersection>96 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>96,-40.5,96,-24</points>
<intersection>-40.5 1</intersection>
<intersection>-24 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>96,-24,139,-24</points>
<connection>
<GID>27</GID>
<name>IN_B_3</name></connection>
<intersection>96 6</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-47.5,113,-47.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108.5,-44.5,113,-44.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-78,276.5,-78</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<connection>
<GID>92</GID>
<name>IN_B_0</name></connection>
<intersection>255 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>255,-78,255,-63</points>
<intersection>-78 1</intersection>
<intersection>-63 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>255,-63,287.5,-63</points>
<connection>
<GID>86</GID>
<name>IN_B_0</name></connection>
<intersection>255 6</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-37,80,-37</points>
<connection>
<GID>14</GID>
<name>OUT_3</name></connection>
<connection>
<GID>22</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-34,80,-34</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<connection>
<GID>22</GID>
<name>IN_B_0</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-92.5,80,-92.5</points>
<intersection>31 5</intersection>
<intersection>80 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>31,-92.5,31,-85</points>
<connection>
<GID>216</GID>
<name>OUT_3</name></connection>
<intersection>-92.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>80,-92.5,80,-84</points>
<connection>
<GID>217</GID>
<name>IN_3</name></connection>
<intersection>-92.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-92.5,80,-83</points>
<connection>
<GID>217</GID>
<name>IN_2</name></connection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-92.5,80,-92.5</points>
<intersection>31 3</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-92.5,31,-87</points>
<connection>
<GID>216</GID>
<name>OUT_2</name></connection>
<intersection>-92.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-36,69.5,-33.5</points>
<intersection>-36 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-33.5,72,-33.5</points>
<connection>
<GID>14</GID>
<name>IN_B_3</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-36,69.5,-36</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-80,276.5,-80</points>
<connection>
<GID>85</GID>
<name>OUT_2</name></connection>
<connection>
<GID>92</GID>
<name>IN_B_2</name></connection>
<intersection>257 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>257,-80,257,-65</points>
<intersection>-80 1</intersection>
<intersection>-65 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>257,-65,287.5,-65</points>
<connection>
<GID>86</GID>
<name>IN_B_2</name></connection>
<intersection>257 6</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-79,276.5,-79</points>
<connection>
<GID>85</GID>
<name>OUT_1</name></connection>
<connection>
<GID>92</GID>
<name>IN_B_1</name></connection>
<intersection>256 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>256,-79,256,-64</points>
<intersection>-79 1</intersection>
<intersection>-64 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>256,-64,287.5,-64</points>
<connection>
<GID>86</GID>
<name>IN_B_1</name></connection>
<intersection>256 8</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-81,276.5,-81</points>
<connection>
<GID>85</GID>
<name>OUT_3</name></connection>
<connection>
<GID>92</GID>
<name>IN_B_3</name></connection>
<intersection>258.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>258.5,-81,258.5,-66</points>
<intersection>-81 1</intersection>
<intersection>-66 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>258.5,-66,287.5,-66</points>
<connection>
<GID>86</GID>
<name>IN_B_3</name></connection>
<intersection>258.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>276.5,-88,276.5,-88</points>
<connection>
<GID>92</GID>
<name>IN_3</name></connection>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-92.5,80,-82</points>
<connection>
<GID>217</GID>
<name>IN_1</name></connection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-92.5,80,-92.5</points>
<intersection>31 3</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-92.5,31,-89</points>
<connection>
<GID>216</GID>
<name>OUT_1</name></connection>
<intersection>-92.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-92.5,80,-81</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-92.5,80,-92.5</points>
<intersection>31 3</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-92.5,31,-91</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>-92.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-53,80,-41</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-53,80,-53</points>
<intersection>30.5 3</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-53,30.5,-50</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>-53 2</intersection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-51.5,80,-42</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-51.5,80,-51.5</points>
<intersection>30.5 3</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-51.5,30.5,-48</points>
<connection>
<GID>19</GID>
<name>OUT_1</name></connection>
<intersection>-51.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88.5,-73,116.5,-73</points>
<connection>
<GID>55</GID>
<name>IN_B_0</name></connection>
<intersection>88.5 9</intersection>
<intersection>95 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>95,-73,95,-58</points>
<intersection>-73 1</intersection>
<intersection>-58 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>95,-58,139,-58</points>
<connection>
<GID>54</GID>
<name>IN_B_0</name></connection>
<intersection>95 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>88.5,-77.5,88.5,-73</points>
<intersection>-77.5 12</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>88,-77.5,88.5,-77.5</points>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<intersection>88.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91,-75,116.5,-75</points>
<connection>
<GID>55</GID>
<name>IN_B_2</name></connection>
<intersection>91 8</intersection>
<intersection>97 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>97,-75,97,-60</points>
<intersection>-75 1</intersection>
<intersection>-60 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>97,-60,139,-60</points>
<connection>
<GID>54</GID>
<name>IN_B_2</name></connection>
<intersection>97 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>91,-79.5,91,-75</points>
<intersection>-79.5 9</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>88,-79.5,91,-79.5</points>
<connection>
<GID>217</GID>
<name>OUT_2</name></connection>
<intersection>91 8</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,-74,116.5,-74</points>
<connection>
<GID>55</GID>
<name>IN_B_1</name></connection>
<intersection>90 10</intersection>
<intersection>96 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>96,-74,96,-59</points>
<intersection>-74 1</intersection>
<intersection>-59 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>96,-59,139,-59</points>
<connection>
<GID>54</GID>
<name>IN_B_1</name></connection>
<intersection>96 8</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>90,-78.5,90,-74</points>
<intersection>-78.5 14</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>88,-78.5,90,-78.5</points>
<connection>
<GID>217</GID>
<name>OUT_1</name></connection>
<intersection>90 10</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-76,116.5,-76</points>
<connection>
<GID>55</GID>
<name>IN_B_3</name></connection>
<intersection>93.5 8</intersection>
<intersection>98.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>98.5,-76,98.5,-61</points>
<intersection>-76 1</intersection>
<intersection>-61 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>98.5,-61,139,-61</points>
<connection>
<GID>54</GID>
<name>IN_B_3</name></connection>
<intersection>98.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>93.5,-80.5,93.5,-76</points>
<intersection>-80.5 9</intersection>
<intersection>-76 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>88,-80.5,93.5,-80.5</points>
<connection>
<GID>217</GID>
<name>OUT_3</name></connection>
<intersection>93.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>116.5,-83,116.5,-83</points>
<connection>
<GID>55</GID>
<name>IN_3</name></connection>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-50.5,79.5,-43</points>
<intersection>-50.5 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-50.5,79.5,-50.5</points>
<intersection>30.5 3</intersection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79.5,-43,80,-43</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>79.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-50.5,30.5,-46</points>
<connection>
<GID>19</GID>
<name>OUT_2</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-49.5,80,-49.5</points>
<intersection>30.5 3</intersection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-49.5,80,-44</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-49.5,30.5,-44</points>
<connection>
<GID>19</GID>
<name>OUT_3</name></connection>
<intersection>-49.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>166.5,-75.5,166.5,-75.5</points>
<connection>
<GID>63</GID>
<name>N_in2</name></connection>
<connection>
<GID>81</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>166.5,-77.5,166.5,-77.5</points>
<connection>
<GID>81</GID>
<name>N_in2</name></connection>
<connection>
<GID>129</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-32.5,72,-32.5</points>
<connection>
<GID>14</GID>
<name>IN_B_2</name></connection>
<intersection>69 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>69,-32.5,69,-32</points>
<connection>
<GID>199</GID>
<name>OUT</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-84.5,214.5,-84</points>
<intersection>-84.5 5</intersection>
<intersection>-84 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>193,-84,214.5,-84</points>
<connection>
<GID>84</GID>
<name>OUT_3</name></connection>
<intersection>214.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>214.5,-84.5,236,-84.5</points>
<connection>
<GID>85</GID>
<name>IN_3</name></connection>
<intersection>214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-86,214.5,-83.5</points>
<intersection>-86 3</intersection>
<intersection>-83.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>193,-86,214.5,-86</points>
<connection>
<GID>84</GID>
<name>OUT_2</name></connection>
<intersection>214.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>214.5,-83.5,236,-83.5</points>
<connection>
<GID>85</GID>
<name>IN_2</name></connection>
<intersection>214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-88,214.5,-82.5</points>
<intersection>-88 3</intersection>
<intersection>-82.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>193,-88,214.5,-88</points>
<connection>
<GID>84</GID>
<name>OUT_1</name></connection>
<intersection>214.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>214.5,-82.5,236,-82.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-71,83,-47</points>
<connection>
<GID>22</GID>
<name>carry_out</name></connection>
<connection>
<GID>217</GID>
<name>carry_in</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-53.5,123.5,-53.5</points>
<intersection>83 0</intersection>
<intersection>123.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123.5,-53.5,123.5,-50.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>-53.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-90,214.5,-81.5</points>
<intersection>-90 3</intersection>
<intersection>-81.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>193,-90,214.5,-90</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>214.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>214.5,-81.5,236,-81.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-27.5,162,-24.5</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-27.5,162,-27.5</points>
<connection>
<GID>27</GID>
<name>OUT_3</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-26.5,162,-25.5</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-26.5,162,-26.5</points>
<connection>
<GID>27</GID>
<name>OUT_2</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>162,-26.5,162,-25.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>-25.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>147,-25.5,162,-25.5</points>
<connection>
<GID>27</GID>
<name>OUT_1</name></connection>
<intersection>162 3</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-27.5,162,-24.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-24.5,162,-24.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>289,-94.5,289,-77.5</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>-77.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>286.5,-77.5,289,-77.5</points>
<intersection>286.5 10</intersection>
<intersection>289 2</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>286.5,-77.5,286.5,-71</points>
<intersection>-77.5 8</intersection>
<intersection>-72 12</intersection>
<intersection>-71 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>286.5,-71,287.5,-71</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>286.5 10</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>286.5,-72,287.5,-72</points>
<connection>
<GID>86</GID>
<name>IN_2</name></connection>
<intersection>286.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>119,-51,121.5,-51</points>
<intersection>119 6</intersection>
<intersection>121.5 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>119,-51,119,-50.5</points>
<connection>
<GID>37</GID>
<name>A_less_B</name></connection>
<intersection>-51 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>121.5,-51,121.5,-50.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>-51 2</intersection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-71.5,239,-52</points>
<connection>
<GID>66</GID>
<name>carry_out</name></connection>
<connection>
<GID>85</GID>
<name>carry_in</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,-58,284.5,-58</points>
<intersection>239 0</intersection>
<intersection>284.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>284.5,-58,284.5,-56</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>-58 1</intersection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295,-32.5,295,-29</points>
<intersection>-32.5 1</intersection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293,-32.5,295,-32.5</points>
<connection>
<GID>67</GID>
<name>OUT_3</name></connection>
<intersection>295 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295,-29,299,-29</points>
<connection>
<GID>114</GID>
<name>IN_3</name></connection>
<intersection>295 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-64.5,163.5,-61.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-61.5,163.5,-61.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-63.5,146.5,-62.5</points>
<intersection>-63.5 1</intersection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>146.5,-63.5,163.5,-63.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>146.5,-62.5,147,-62.5</points>
<connection>
<GID>54</GID>
<name>OUT_1</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-63.5,163.5,-62.5</points>
<connection>
<GID>73</GID>
<name>IN_2</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-63.5,163.5,-63.5</points>
<connection>
<GID>54</GID>
<name>OUT_2</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164,-64.5,164,-61.5</points>
<intersection>-64.5 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-64.5,164,-64.5</points>
<connection>
<GID>54</GID>
<name>OUT_3</name></connection>
<intersection>164 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163.5,-61.5,164,-61.5</points>
<connection>
<GID>73</GID>
<name>IN_3</name></connection>
<intersection>164 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-88.5,122.5,-86</points>
<connection>
<GID>55</GID>
<name>A_less_B</name></connection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-88.5,123,-88.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166,-79.5,166.5,-79.5</points>
<connection>
<GID>174</GID>
<name>N_in3</name></connection>
<connection>
<GID>129</GID>
<name>N_in2</name></connection>
<intersection>166 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>166,-79.5,166,-78.5</points>
<intersection>-79.5 1</intersection>
<intersection>-78.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>165.5,-78.5,166,-78.5</points>
<connection>
<GID>129</GID>
<name>N_in0</name></connection>
<intersection>166 4</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-55,142,-34</points>
<connection>
<GID>54</GID>
<name>carry_in</name></connection>
<connection>
<GID>27</GID>
<name>carry_out</name></connection>
<intersection>-54.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>104,-54.5,142,-54.5</points>
<intersection>104 9</intersection>
<intersection>142 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>104,-81,104,-54.5</points>
<intersection>-81 10</intersection>
<intersection>-54.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>104,-81,109,-81</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>104 9</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295,-31.5,295,-30</points>
<intersection>-31.5 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293,-31.5,295,-31.5</points>
<connection>
<GID>67</GID>
<name>OUT_2</name></connection>
<intersection>295 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295,-30,299,-30</points>
<connection>
<GID>114</GID>
<name>IN_2</name></connection>
<intersection>295 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-79,109,-79</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>293,-31,299,-31</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>293 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>293,-31,293,-30.5</points>
<connection>
<GID>67</GID>
<name>OUT_1</name></connection>
<intersection>-31 1</intersection></vsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296,-32,296,-29.5</points>
<intersection>-32 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293,-29.5,296,-29.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>296 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>296,-32,299,-32</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>296 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>279,-56,282.5,-56</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>279 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>279,-56,279,-55.5</points>
<connection>
<GID>75</GID>
<name>A_less_B</name></connection>
<intersection>-56 2</intersection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>115,-80,116.5,-80</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>78</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-69.5,298,-66.5</points>
<intersection>-69.5 2</intersection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-66.5,298,-66.5</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>298 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>298,-69.5,300.5,-69.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>298 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-68.5,298,-67.5</points>
<intersection>-68.5 1</intersection>
<intersection>-67.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>298,-68.5,300.5,-68.5</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>298 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295.5,-67.5,298,-67.5</points>
<connection>
<GID>86</GID>
<name>OUT_1</name></connection>
<intersection>298 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-68.5,298,-67.5</points>
<intersection>-68.5 1</intersection>
<intersection>-67.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-68.5,298,-68.5</points>
<connection>
<GID>86</GID>
<name>OUT_2</name></connection>
<intersection>298 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>298,-67.5,300.5,-67.5</points>
<connection>
<GID>120</GID>
<name>IN_2</name></connection>
<intersection>298 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-69.5,298,-66.5</points>
<intersection>-69.5 1</intersection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-69.5,298,-69.5</points>
<connection>
<GID>86</GID>
<name>OUT_3</name></connection>
<intersection>298 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>298,-66.5,300.5,-66.5</points>
<connection>
<GID>120</GID>
<name>IN_3</name></connection>
<intersection>298 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282.5,-93.5,282.5,-91</points>
<connection>
<GID>92</GID>
<name>A_less_B</name></connection>
<intersection>-93.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282.5,-93.5,283,-93.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>282.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-95.5,239,-87.5</points>
<connection>
<GID>85</GID>
<name>carry_out</name></connection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,-95.5,283,-95.5</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-60,288,-39</points>
<connection>
<GID>67</GID>
<name>carry_out</name></connection>
<intersection>-60 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>264,-60,290.5,-60</points>
<connection>
<GID>86</GID>
<name>carry_in</name></connection>
<intersection>264 6</intersection>
<intersection>288 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>264,-86,264,-60</points>
<intersection>-86 7</intersection>
<intersection>-60 3</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>264,-86,269,-86</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>264 6</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>269,-84,269,-84</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>275,-85,276.5,-85</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-73.5,172,-9.5</points>
<intersection>-73.5 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-9.5,172,-9.5</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>172 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,-73.5,172,-73.5</points>
<connection>
<GID>63</GID>
<name>N_in3</name></connection>
<intersection>172 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-44.5,122.5,-32</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>-36 21</intersection>
<intersection>-32 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>122.5,-32,131.5,-32</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>122.5,-36,131.5,-36</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-35,138.5,-30</points>
<intersection>-35 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-30,139,-30</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-35,138.5,-35</points>
<connection>
<GID>191</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-31,138,-29</points>
<intersection>-31 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-29,139,-29</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-31,138,-31</points>
<connection>
<GID>190</GID>
<name>OUT</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-28,138,-27</points>
<intersection>-28 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-28,139,-28</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-27,138,-27</points>
<connection>
<GID>189</GID>
<name>OUT</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-39,139,-31</points>
<connection>
<GID>27</GID>
<name>IN_3</name></connection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-39,139,-39</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-31.5,69.5,-28</points>
<intersection>-31.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-31.5,72,-31.5</points>
<connection>
<GID>14</GID>
<name>IN_B_1</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-28,69.5,-28</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-28,131.5,-28</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-40,131.5,-40</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-89.5,129,-68</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>-72 21</intersection>
<intersection>-68 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>129,-68,132,-68</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>129,-72,132,-72</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-64,132,-64</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<connection>
<GID>210</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-76,132,-76</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<connection>
<GID>213</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-30.5,69.5,-24</points>
<intersection>-30.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-24,69.5,-24</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-30.5,72,-30.5</points>
<connection>
<GID>14</GID>
<name>IN_B_0</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-80.5,62,-15</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>-80.5 136</intersection>
<intersection>-40.5 31</intersection>
<intersection>-35 101</intersection>
<intersection>-31 39</intersection>
<intersection>-27 29</intersection>
<intersection>-23 28</intersection>
<intersection>-15 30</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>62,-23,63,-23</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>62,-27,63,-27</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>62,-15,142,-15</points>
<intersection>62 0</intersection>
<intersection>127.5 37</intersection>
<intersection>142 226</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>62,-40.5,75,-40.5</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<intersection>62 0</intersection>
<intersection>70.5 224</intersection>
<intersection>75 222</intersection></hsegment>
<vsegment>
<ID>37</ID>
<points>127.5,-74,127.5,-15</points>
<intersection>-74 90</intersection>
<intersection>-70 98</intersection>
<intersection>-66 95</intersection>
<intersection>-62 96</intersection>
<intersection>-38 40</intersection>
<intersection>-34 48</intersection>
<intersection>-30 45</intersection>
<intersection>-26 228</intersection>
<intersection>-15 30</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>62,-31,63,-31</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>127.5,-38,131.5,-38</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>127.5,-30,131.5,-30</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>127.5,-34,131.5,-34</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>90</ID>
<points>127.5,-74,132,-74</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>95</ID>
<points>127.5,-66,132,-66</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>96</ID>
<points>127.5,-62,132,-62</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>98</ID>
<points>127.5,-70,132,-70</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment>
<hsegment>
<ID>101</ID>
<points>62,-35,63,-35</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>136</ID>
<points>62,-80.5,72,-80.5</points>
<connection>
<GID>41</GID>
<name>IN_3</name></connection>
<intersection>62 0</intersection>
<intersection>71.5 218</intersection></hsegment>
<vsegment>
<ID>218</ID>
<points>71.5,-80.5,71.5,-77.5</points>
<intersection>-80.5 136</intersection>
<intersection>-77.5 221</intersection></vsegment>
<hsegment>
<ID>221</ID>
<points>71.5,-77.5,75,-77.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>71.5 218</intersection>
<intersection>75 223</intersection></hsegment>
<vsegment>
<ID>222</ID>
<points>75,-40.5,75,-27.5</points>
<connection>
<GID>14</GID>
<name>carry_in</name></connection>
<intersection>-40.5 31</intersection></vsegment>
<vsegment>
<ID>223</ID>
<points>75,-77.5,75,-67.5</points>
<connection>
<GID>41</GID>
<name>carry_in</name></connection>
<intersection>-77.5 221</intersection></vsegment>
<vsegment>
<ID>224</ID>
<points>70.5,-40.5,70.5,-37.5</points>
<intersection>-40.5 31</intersection>
<intersection>-37.5 225</intersection></vsegment>
<hsegment>
<ID>225</ID>
<points>70.5,-37.5,72,-37.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>70.5 224</intersection></hsegment>
<vsegment>
<ID>226</ID>
<points>142,-18,142,-15</points>
<connection>
<GID>27</GID>
<name>carry_in</name></connection>
<intersection>-15 30</intersection></vsegment>
<hsegment>
<ID>228</ID>
<points>127.5,-26,131.5,-26</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>127.5 37</intersection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>518,-18,518,33</points>
<connection>
<GID>672</GID>
<name>OUT_0</name></connection>
<intersection>3 9</intersection>
<intersection>16.5 4</intersection>
<intersection>33 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>511,16.5,518,16.5</points>
<intersection>511 7</intersection>
<intersection>518 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>512,33,518,33</points>
<intersection>512 8</intersection>
<intersection>517.5 13</intersection>
<intersection>518 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>511,15,511,19</points>
<connection>
<GID>313</GID>
<name>load</name></connection>
<intersection>16.5 4</intersection>
<intersection>19 16</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>512,32,512,33</points>
<connection>
<GID>312</GID>
<name>load</name></connection>
<intersection>33 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>510,3,518,3</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>511 11</intersection>
<intersection>518 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>511,-1,511,3</points>
<connection>
<GID>325</GID>
<name>load</name></connection>
<intersection>3 9</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>517.5,33,517.5,37.5</points>
<intersection>33 6</intersection>
<intersection>37.5 20</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>509.5,19,511,19</points>
<intersection>509.5 21</intersection>
<intersection>511 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>510,37.5,517.5,37.5</points>
<intersection>510 22</intersection>
<intersection>517.5 13</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>509.5,19,509.5,20</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>19 16</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>510,37,510,37.5</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>37.5 20</intersection></vsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-76,80,-76</points>
<connection>
<GID>41</GID>
<name>OUT_2</name></connection>
<connection>
<GID>217</GID>
<name>IN_B_2</name></connection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-74,80,-74</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<connection>
<GID>217</GID>
<name>IN_B_0</name></connection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-75,80,-75</points>
<connection>
<GID>41</GID>
<name>OUT_1</name></connection>
<connection>
<GID>217</GID>
<name>IN_B_1</name></connection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-75,139,-68</points>
<connection>
<GID>54</GID>
<name>IN_3</name></connection>
<intersection>-75 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138,-75,139,-75</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-77,80,-77</points>
<connection>
<GID>41</GID>
<name>OUT_3</name></connection>
<connection>
<GID>217</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-65,138.5,-63</points>
<intersection>-65 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-65,139,-65</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-63,138.5,-63</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-67,138,-66</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-66,139,-66</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-71,138.5,-67</points>
<intersection>-71 4</intersection>
<intersection>-67 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>138.5,-67,139,-67</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>138,-71,138.5,-71</points>
<connection>
<GID>212</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-37,61,-30.5</points>
<intersection>-37 5</intersection>
<intersection>-30.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>57,-30.5,61,-30.5</points>
<connection>
<GID>17</GID>
<name>OUT_3</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61,-37,63,-37</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-33,61,-32.5</points>
<intersection>-33 5</intersection>
<intersection>-32.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>57,-32.5,61,-32.5</points>
<connection>
<GID>17</GID>
<name>OUT_2</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61,-33,63,-33</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-34.5,61,-29</points>
<intersection>-34.5 4</intersection>
<intersection>-29 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>57,-34.5,61,-34.5</points>
<connection>
<GID>17</GID>
<name>OUT_1</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61,-29,63,-29</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-36.5,61,-25</points>
<intersection>-36.5 4</intersection>
<intersection>-25 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>57,-36.5,61,-36.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61,-25,63,-25</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-70.5,70,-65</points>
<intersection>-70.5 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-70.5,72,-70.5</points>
<connection>
<GID>41</GID>
<name>IN_B_0</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-65,70,-65</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393.5,-11.5,393.5,-4</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<intersection>-11.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>384.5,-11.5,393.5,-11.5</points>
<connection>
<GID>228</GID>
<name>IN_B_0</name></connection>
<intersection>393.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>383.5,-11.5,383.5,-7.5</points>
<connection>
<GID>228</GID>
<name>IN_B_1</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>389.5,-7.5,389.5,-4</points>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>383.5,-7.5,389.5,-7.5</points>
<intersection>383.5 0</intersection>
<intersection>389.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>382.5,-11.5,382.5,-4</points>
<connection>
<GID>228</GID>
<name>IN_B_2</name></connection>
<intersection>-4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>382.5,-4,385.5,-4</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<intersection>382.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-71.5,69.5,-69</points>
<intersection>-71.5 2</intersection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-69,69.5,-69</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-71.5,72,-71.5</points>
<connection>
<GID>41</GID>
<name>IN_B_1</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381.5,-11.5,381.5,-4</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<connection>
<GID>228</GID>
<name>IN_B_3</name></connection></vsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-73,70,-72.5</points>
<intersection>-73 1</intersection>
<intersection>-72.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-73,70,-73</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-72.5,72,-72.5</points>
<connection>
<GID>41</GID>
<name>IN_B_2</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-77,70,-73.5</points>
<intersection>-77 1</intersection>
<intersection>-73.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-77,70,-77</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-73.5,72,-73.5</points>
<connection>
<GID>41</GID>
<name>IN_B_3</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-10.5,-106.5,-10</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-106.5,-10,-88.5,-10</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-104.5,-12,-104.5,-10.5</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-104.5,-12,-88.5,-12</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>-104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79.5,-39,-54.5,-39</points>
<connection>
<GID>252</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<intersection>-75 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-75,-39,-75,-22.5</points>
<intersection>-39 1</intersection>
<intersection>-22.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-75,-22.5,-28.5,-22.5</points>
<connection>
<GID>242</GID>
<name>IN_B_0</name></connection>
<intersection>-75 6</intersection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-78,60,-71.5</points>
<intersection>-78 3</intersection>
<intersection>-71.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>60,-78,62,-78</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>55.5,-71.5,60,-71.5</points>
<connection>
<GID>214</GID>
<name>OUT_3</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-74,60,-73.5</points>
<intersection>-74 3</intersection>
<intersection>-73.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>60,-74,62,-74</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>55.5,-73.5,60,-73.5</points>
<connection>
<GID>214</GID>
<name>OUT_2</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-75.5,60,-70</points>
<intersection>-75.5 4</intersection>
<intersection>-70 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>60,-70,62,-70</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>55.5,-75.5,60,-75.5</points>
<connection>
<GID>214</GID>
<name>OUT_1</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-77.5,60,-66</points>
<intersection>-77.5 4</intersection>
<intersection>-66 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>60,-66,62,-66</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>55.5,-77.5,60,-77.5</points>
<connection>
<GID>214</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>343,4.5,402.5,4.5</points>
<intersection>343 18</intersection>
<intersection>345 21</intersection>
<intersection>351 25</intersection>
<intersection>355 24</intersection>
<intersection>359 23</intersection>
<intersection>363 22</intersection>
<intersection>374.5 5</intersection>
<intersection>376.5 8</intersection>
<intersection>382.5 26</intersection>
<intersection>386.5 27</intersection>
<intersection>390.5 28</intersection>
<intersection>394.5 29</intersection>
<intersection>402.5 9</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>374.5,-11.5,374.5,4.5</points>
<connection>
<GID>228</GID>
<name>IN_3</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>376.5,-11.5,376.5,4.5</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>402.5,4.5,402.5,36.5</points>
<intersection>4.5 1</intersection>
<intersection>36.5 11</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>365.5,36.5,365.5,37.5</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>36.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>363,36.5,402.5,36.5</points>
<connection>
<GID>259</GID>
<name>nQ</name></connection>
<intersection>365.5 10</intersection>
<intersection>402.5 9</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>343,-11.5,343,4.5</points>
<connection>
<GID>282</GID>
<name>IN_3</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>345,-11.5,345,4.5</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>363,2,363,4.5</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>359,2,359,4.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>355,2,355,4.5</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>351,2,351,4.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>382.5,2,382.5,4.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>386.5,2,386.5,4.5</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>390.5,2,390.5,4.5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>394.5,2,394.5,4.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>4.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79.5,-41,-54.5,-41</points>
<connection>
<GID>252</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>236</GID>
<name>OUT_2</name></connection>
<intersection>-73 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-73,-41,-73,-24.5</points>
<intersection>-41 1</intersection>
<intersection>-24.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-73,-24.5,-28.5,-24.5</points>
<connection>
<GID>242</GID>
<name>IN_B_2</name></connection>
<intersection>-73 6</intersection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79.5,-40,-54.5,-40</points>
<connection>
<GID>252</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>236</GID>
<name>OUT_1</name></connection>
<intersection>-74 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-74,-40,-74,-23.5</points>
<intersection>-40 1</intersection>
<intersection>-23.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-74,-23.5,-28.5,-23.5</points>
<connection>
<GID>242</GID>
<name>IN_B_1</name></connection>
<intersection>-74 8</intersection></hsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379,-22,379,-19.5</points>
<connection>
<GID>228</GID>
<name>OUT_2</name></connection>
<intersection>-22 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>373.5,-22,379,-22</points>
<intersection>373.5 16</intersection>
<intersection>379 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>373.5,-25,373.5,-22</points>
<connection>
<GID>241</GID>
<name>IN_B_2</name></connection>
<intersection>-22 5</intersection></vsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-90.5,83,-87</points>
<connection>
<GID>217</GID>
<name>carry_out</name></connection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-90.5,123,-90.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381,-25,381,-19.5</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>-25 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>375.5,-25,381,-25</points>
<connection>
<GID>241</GID>
<name>IN_B_0</name></connection>
<intersection>381 0</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372.5,-25,372.5,-19.5</points>
<connection>
<GID>241</GID>
<name>IN_B_3</name></connection>
<intersection>-19.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>372.5,-19.5,378,-19.5</points>
<connection>
<GID>228</GID>
<name>OUT_3</name></connection>
<intersection>372.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,-23,380,-19.5</points>
<connection>
<GID>228</GID>
<name>OUT_1</name></connection>
<intersection>-23 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>374.5,-23,380,-23</points>
<intersection>374.5 16</intersection>
<intersection>380 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>374.5,-25,374.5,-23</points>
<connection>
<GID>241</GID>
<name>IN_B_1</name></connection>
<intersection>-23 5</intersection></vsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79.5,-42,-54.5,-42</points>
<connection>
<GID>252</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>236</GID>
<name>OUT_3</name></connection>
<intersection>-71.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-71.5,-42,-71.5,-25.5</points>
<intersection>-42 1</intersection>
<intersection>-25.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-71.5,-25.5,-28.5,-25.5</points>
<connection>
<GID>242</GID>
<name>IN_B_3</name></connection>
<intersection>-71.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-49,-54.5,-49</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<connection>
<GID>252</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59,-46,-54.5,-46</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<connection>
<GID>252</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>523.5,-27,523.5,22</points>
<intersection>-27 16</intersection>
<intersection>-23 4</intersection>
<intersection>5 3</intersection>
<intersection>22 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>511,5,523.5,5</points>
<connection>
<GID>313</GID>
<name>clock</name></connection>
<intersection>523.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>495.5,-23,523.5,-23</points>
<connection>
<GID>670</GID>
<name>CLK</name></connection>
<intersection>511 7</intersection>
<intersection>523.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>512,22,523.5,22</points>
<connection>
<GID>312</GID>
<name>clock</name></connection>
<intersection>523.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>511,-23,511,-11</points>
<connection>
<GID>325</GID>
<name>clock</name></connection>
<intersection>-23 4</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>523.5,-27,533,-27</points>
<connection>
<GID>311</GID>
<name>clock</name></connection>
<intersection>523.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>508.5,-1,508.5,5</points>
<connection>
<GID>325</GID>
<name>carry_in</name></connection>
<connection>
<GID>313</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,21.5,366.5,40.5</points>
<connection>
<GID>264</GID>
<name>N_in2</name></connection>
<intersection>26.5 12</intersection>
<intersection>37.5 13</intersection>
<intersection>40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>363,40.5,366.5,40.5</points>
<connection>
<GID>259</GID>
<name>Q</name></connection>
<intersection>366.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>366.5,26.5,367.5,26.5</points>
<connection>
<GID>266</GID>
<name>N_in1</name></connection>
<intersection>366.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>366.5,37.5,367.5,37.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>366.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>357,36.5,357,40.5</points>
<connection>
<GID>259</GID>
<name>clock</name></connection>
<connection>
<GID>259</GID>
<name>K</name></connection>
<connection>
<GID>259</GID>
<name>J</name></connection>
<connection>
<GID>257</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,24.5,366.5,31.5</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>365.5,24.5,369.5,24.5</points>
<connection>
<GID>268</GID>
<name>N_in1</name></connection>
<connection>
<GID>261</GID>
<name>N_in1</name></connection>
<connection>
<GID>272</GID>
<name>N_in1</name></connection>
<intersection>366.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-136.5,-94,-87.5,-94</points>
<intersection>-136.5 5</intersection>
<intersection>-87.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-136.5,-94,-136.5,-86.5</points>
<connection>
<GID>238</GID>
<name>OUT_3</name></connection>
<intersection>-94 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-87.5,-94,-87.5,-85.5</points>
<connection>
<GID>240</GID>
<name>IN_3</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-94,-87.5,-84.5</points>
<connection>
<GID>240</GID>
<name>IN_2</name></connection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-136.5,-94,-87.5,-94</points>
<intersection>-136.5 3</intersection>
<intersection>-87.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-136.5,-94,-136.5,-88.5</points>
<connection>
<GID>238</GID>
<name>OUT_2</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362,-11.5,362,-4</points>
<connection>
<GID>281</GID>
<name>OUT</name></connection>
<intersection>-11.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>353,-11.5,362,-11.5</points>
<connection>
<GID>282</GID>
<name>IN_B_0</name></connection>
<intersection>362 0</intersection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-11.5,352,-7.5</points>
<connection>
<GID>282</GID>
<name>IN_B_1</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>358,-7.5,358,-4</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>352,-7.5,358,-7.5</points>
<intersection>352 0</intersection>
<intersection>358 1</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351,-11.5,351,-4</points>
<connection>
<GID>282</GID>
<name>IN_B_2</name></connection>
<intersection>-4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>351,-4,354,-4</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<intersection>351 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-11.5,350,-4</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<connection>
<GID>282</GID>
<name>IN_B_3</name></connection></vsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520.5,-13,520.5,-7.5</points>
<intersection>-13 3</intersection>
<intersection>-7.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>520.5,-13,528,-13</points>
<connection>
<GID>410</GID>
<name>IN_1</name></connection>
<intersection>520.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>513.5,-7.5,520.5,-7.5</points>
<connection>
<GID>325</GID>
<name>OUT_3</name></connection>
<intersection>520.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347.5,-22,347.5,-19.5</points>
<connection>
<GID>282</GID>
<name>OUT_2</name></connection>
<intersection>-22 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>342,-22,347.5,-22</points>
<intersection>342 12</intersection>
<intersection>347.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>342,-25,342,-22</points>
<connection>
<GID>283</GID>
<name>IN_B_2</name></connection>
<intersection>-22 5</intersection></vsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,-23,349.5,-19.5</points>
<connection>
<GID>282</GID>
<name>OUT_0</name></connection>
<intersection>-23 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>344,-23,349.5,-23</points>
<intersection>344 9</intersection>
<intersection>349.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>344,-25,344,-23</points>
<connection>
<GID>283</GID>
<name>IN_B_0</name></connection>
<intersection>-23 5</intersection></vsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341,-25,341,-21.5</points>
<connection>
<GID>283</GID>
<name>IN_B_3</name></connection>
<intersection>-21.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>341,-21.5,346.5,-21.5</points>
<intersection>341 0</intersection>
<intersection>346.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>346.5,-21.5,346.5,-19.5</points>
<connection>
<GID>282</GID>
<name>OUT_3</name></connection>
<intersection>-21.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>348.5,-22.5,348.5,-19.5</points>
<connection>
<GID>282</GID>
<name>OUT_1</name></connection>
<intersection>-22.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>343,-22.5,348.5,-22.5</points>
<intersection>343 6</intersection>
<intersection>348.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>343,-25,343,-22.5</points>
<connection>
<GID>283</GID>
<name>IN_B_1</name></connection>
<intersection>-22.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-94,-87.5,-83.5</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-136.5,-94,-87.5,-94</points>
<intersection>-136.5 3</intersection>
<intersection>-87.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-136.5,-94,-136.5,-90.5</points>
<connection>
<GID>238</GID>
<name>OUT_1</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-94,-87.5,-82.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-136.5,-94,-87.5,-94</points>
<intersection>-136.5 3</intersection>
<intersection>-87.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-136.5,-94,-136.5,-92.5</points>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349,2,349,13.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>13.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>349,13.5,384,13.5</points>
<intersection>349 0</intersection>
<intersection>384 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>384,13.5,384,27.5</points>
<intersection>13.5 2</intersection>
<intersection>27.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>381.5,27.5,384,27.5</points>
<connection>
<GID>246</GID>
<name>OUT_3</name></connection>
<intersection>384 3</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>353,12.5,383.5,12.5</points>
<intersection>353 4</intersection>
<intersection>383.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383.5,12.5,383.5,25.5</points>
<intersection>12.5 1</intersection>
<intersection>25.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>381.5,25.5,383.5,25.5</points>
<connection>
<GID>246</GID>
<name>OUT_2</name></connection>
<intersection>383.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>353,2,353,12.5</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,2,357,11.5</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,11.5,383,11.5</points>
<intersection>357 0</intersection>
<intersection>383 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383,11.5,383,23.5</points>
<intersection>11.5 1</intersection>
<intersection>23.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>381.5,23.5,383,23.5</points>
<connection>
<GID>246</GID>
<name>OUT_1</name></connection>
<intersection>383 2</intersection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361,2,361,10.5</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361,10.5,381.5,10.5</points>
<intersection>361 0</intersection>
<intersection>381.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>381.5,10.5,381.5,21.5</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380.5,2,380.5,9</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380.5,9,400.5,9</points>
<intersection>380.5 0</intersection>
<intersection>400.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>400.5,9,400.5,27</points>
<intersection>9 1</intersection>
<intersection>27 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>396,27,400.5,27</points>
<connection>
<GID>248</GID>
<name>OUT_3</name></connection>
<intersection>400.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384.5,2,384.5,8.5</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384.5,8.5,399.5,8.5</points>
<intersection>384.5 0</intersection>
<intersection>399.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>399.5,8.5,399.5,25</points>
<intersection>8.5 1</intersection>
<intersection>25 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>396,25,399.5,25</points>
<connection>
<GID>248</GID>
<name>OUT_2</name></connection>
<intersection>399.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>388.5,2,388.5,7.5</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>388.5,7.5,398.5,7.5</points>
<intersection>388.5 0</intersection>
<intersection>398.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>398.5,7.5,398.5,23</points>
<intersection>7.5 1</intersection>
<intersection>23 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>396,23,398.5,23</points>
<connection>
<GID>248</GID>
<name>OUT_1</name></connection>
<intersection>398.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>392.5,2,392.5,7</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>392.5,7,397.5,7</points>
<intersection>392.5 0</intersection>
<intersection>397.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>397.5,7,397.5,21</points>
<intersection>7 1</intersection>
<intersection>21 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>396,21,397.5,21</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>397.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361.5,15.5,361.5,27.5</points>
<intersection>15.5 2</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360.5,27.5,361.5,27.5</points>
<connection>
<GID>245</GID>
<name>OUT_3</name></connection>
<intersection>361.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>361.5,15.5,365.5,15.5</points>
<intersection>361.5 0</intersection>
<intersection>365.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>365.5,-25,365.5,15.5</points>
<connection>
<GID>241</GID>
<name>IN_3</name></connection>
<intersection>15.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,-25,366.5,16</points>
<connection>
<GID>241</GID>
<name>IN_2</name></connection>
<intersection>16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>362.5,16,366.5,16</points>
<intersection>362.5 2</intersection>
<intersection>366.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>362.5,16,362.5,25.5</points>
<intersection>16 1</intersection>
<intersection>25.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>360.5,25.5,362.5,25.5</points>
<connection>
<GID>245</GID>
<name>OUT_2</name></connection>
<intersection>362.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363,16.5,363,23.5</points>
<intersection>16.5 2</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360.5,23.5,363,23.5</points>
<connection>
<GID>245</GID>
<name>OUT_1</name></connection>
<intersection>363 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>363,16.5,367.5,16.5</points>
<intersection>363 0</intersection>
<intersection>367.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>367.5,-25,367.5,16.5</points>
<connection>
<GID>241</GID>
<name>IN_1</name></connection>
<intersection>16.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363.5,17,363.5,21.5</points>
<intersection>17 2</intersection>
<intersection>21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360.5,21.5,363.5,21.5</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>363.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>363.5,17,368.5,17</points>
<intersection>363.5 0</intersection>
<intersection>368.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>368.5,-25,368.5,17</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>17 2</intersection></vsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,-25,334,17</points>
<connection>
<GID>283</GID>
<name>IN_3</name></connection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>334,17,350.5,17</points>
<intersection>334 0</intersection>
<intersection>350.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350.5,17,350.5,27.5</points>
<intersection>17 1</intersection>
<intersection>27.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>349,27.5,350.5,27.5</points>
<connection>
<GID>244</GID>
<name>OUT_3</name></connection>
<intersection>350.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335,-25,335,16.5</points>
<connection>
<GID>283</GID>
<name>IN_2</name></connection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>335,16.5,350,16.5</points>
<intersection>335 0</intersection>
<intersection>350 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350,16.5,350,25.5</points>
<intersection>16.5 1</intersection>
<intersection>25.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>349,25.5,350,25.5</points>
<connection>
<GID>244</GID>
<name>OUT_2</name></connection>
<intersection>350 2</intersection></hsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336,-25,336,16</points>
<connection>
<GID>283</GID>
<name>IN_1</name></connection>
<intersection>16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>336,16,349.5,16</points>
<intersection>336 0</intersection>
<intersection>349.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>349.5,16,349.5,23.5</points>
<intersection>16 1</intersection>
<intersection>23.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>349,23.5,349.5,23.5</points>
<connection>
<GID>244</GID>
<name>OUT_1</name></connection>
<intersection>349.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-25,337,15.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>337,15.5,349,15.5</points>
<intersection>337 0</intersection>
<intersection>349 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>349,15.5,349,21.5</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362.5,-40.5,362.5,-35</points>
<connection>
<GID>284</GID>
<name>IN_B_2</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>362.5,-35,370,-35</points>
<intersection>362.5 0</intersection>
<intersection>370 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>370,-49,370,-33</points>
<connection>
<GID>241</GID>
<name>OUT_2</name></connection>
<connection>
<GID>288</GID>
<name>IN_B_2</name></connection>
<intersection>-35 1</intersection></vsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363.5,-40.5,363.5,-36</points>
<connection>
<GID>284</GID>
<name>IN_B_1</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>363.5,-36,371,-36</points>
<intersection>363.5 0</intersection>
<intersection>371 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>371,-49,371,-33</points>
<connection>
<GID>241</GID>
<name>OUT_1</name></connection>
<connection>
<GID>288</GID>
<name>IN_B_1</name></connection>
<intersection>-36 1</intersection></vsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-49,372,-33</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<connection>
<GID>288</GID>
<name>IN_B_0</name></connection>
<intersection>-36.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>364.5,-36.5,372,-36.5</points>
<intersection>364.5 6</intersection>
<intersection>372 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>364.5,-40.5,364.5,-36.5</points>
<connection>
<GID>284</GID>
<name>IN_B_0</name></connection>
<intersection>-36.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361.5,-40.5,361.5,-34.5</points>
<connection>
<GID>284</GID>
<name>IN_B_3</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361.5,-34.5,369,-34.5</points>
<intersection>361.5 0</intersection>
<intersection>369 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>369,-49,369,-33</points>
<connection>
<GID>241</GID>
<name>OUT_3</name></connection>
<connection>
<GID>288</GID>
<name>IN_B_3</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-54.5,-87.5,-42.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-137,-54.5,-87.5,-54.5</points>
<intersection>-137 3</intersection>
<intersection>-87.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-137,-54.5,-137,-51.5</points>
<intersection>-54.5 2</intersection>
<intersection>-51.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-137.5,-51.5,-137,-51.5</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>-137 3</intersection></hsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354.5,-40.5,354.5,-40.5</points>
<connection>
<GID>284</GID>
<name>IN_3</name></connection>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357.5,-40.5,357.5,-40.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-53,-87.5,-43.5</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-137,-53,-87.5,-53</points>
<intersection>-137 3</intersection>
<intersection>-87.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-137,-53,-137,-49.5</points>
<intersection>-53 2</intersection>
<intersection>-49.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-137.5,-49.5,-137,-49.5</points>
<connection>
<GID>232</GID>
<name>OUT_1</name></connection>
<intersection>-137 3</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331,-40,331,-34.5</points>
<connection>
<GID>290</GID>
<name>IN_B_2</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>331,-34.5,338.5,-34.5</points>
<intersection>331 0</intersection>
<intersection>338.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>338.5,-49,338.5,-33</points>
<connection>
<GID>283</GID>
<name>OUT_2</name></connection>
<connection>
<GID>297</GID>
<name>IN_B_2</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,-40,332,-35.5</points>
<connection>
<GID>290</GID>
<name>IN_B_1</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>332,-35.5,339.5,-35.5</points>
<intersection>332 0</intersection>
<intersection>339.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>339.5,-49,339.5,-33</points>
<connection>
<GID>283</GID>
<name>OUT_1</name></connection>
<connection>
<GID>297</GID>
<name>IN_B_1</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>340.5,-49,340.5,-33</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<connection>
<GID>297</GID>
<name>IN_B_0</name></connection>
<intersection>-36 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>333,-36,340.5,-36</points>
<intersection>333 6</intersection>
<intersection>340.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>333,-40,333,-36</points>
<connection>
<GID>290</GID>
<name>IN_B_0</name></connection>
<intersection>-36 4</intersection></vsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,-40,330,-34</points>
<connection>
<GID>290</GID>
<name>IN_B_3</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>330,-34,337.5,-34</points>
<intersection>330 0</intersection>
<intersection>337.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>337.5,-49,337.5,-33</points>
<connection>
<GID>283</GID>
<name>OUT_3</name></connection>
<connection>
<GID>297</GID>
<name>IN_B_3</name></connection>
<intersection>-34 1</intersection></vsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323,-40,323,-40</points>
<connection>
<GID>290</GID>
<name>IN_3</name></connection>
<connection>
<GID>295</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520.5,-9,520.5,-6.5</points>
<intersection>-9 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,-6.5,520.5,-6.5</points>
<connection>
<GID>325</GID>
<name>OUT_2</name></connection>
<intersection>520.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>520.5,-9,528,-9</points>
<connection>
<GID>409</GID>
<name>IN_1</name></connection>
<intersection>520.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520.5,-5.5,520.5,-5</points>
<intersection>-5.5 1</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,-5.5,520.5,-5.5</points>
<connection>
<GID>325</GID>
<name>OUT_1</name></connection>
<intersection>520.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>520.5,-5,528,-5</points>
<connection>
<GID>408</GID>
<name>IN_1</name></connection>
<intersection>520.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>314.5,-48,332.5,-48</points>
<intersection>314.5 8</intersection>
<intersection>320 3</intersection>
<intersection>331.5 13</intersection>
<intersection>332.5 14</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>320,-48,320,-46</points>
<connection>
<GID>290</GID>
<name>A_less_B</name></connection>
<intersection>-48 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>314.5,-52.5,314.5,-48</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>-48 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>331.5,-49,331.5,-48</points>
<connection>
<GID>297</GID>
<name>IN_2</name></connection>
<intersection>-48 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>332.5,-49,332.5,-48</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>-48 1</intersection></vsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>349,-58.5,372.5,-58.5</points>
<connection>
<GID>307</GID>
<name>OUT_0</name></connection>
<intersection>349 26</intersection>
<intersection>360.5 39</intersection>
<intersection>364.5 27</intersection>
<intersection>368.5 28</intersection>
<intersection>372.5 29</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>349,-69,349,-58.5</points>
<intersection>-69 30</intersection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>364.5,-60,364.5,-58.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>368.5,-60,368.5,-58.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>372.5,-60,372.5,-58.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>349,-69,357.5,-69</points>
<intersection>349 26</intersection>
<intersection>355.5 42</intersection>
<intersection>357.5 32</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>357.5,-70,357.5,-69</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>-69 30</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>360.5,-60,360.5,-58.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>355.5,-70,355.5,-69</points>
<connection>
<GID>302</GID>
<name>IN_3</name></connection>
<intersection>-69 30</intersection></vsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,-74.5,-51,-74.5</points>
<connection>
<GID>275</GID>
<name>IN_B_0</name></connection>
<intersection>-79 9</intersection>
<intersection>-72.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-72.5,-74.5,-72.5,-59.5</points>
<intersection>-74.5 1</intersection>
<intersection>-59.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-72.5,-59.5,-28.5,-59.5</points>
<connection>
<GID>273</GID>
<name>IN_B_0</name></connection>
<intersection>-72.5 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-79,-79,-79,-74.5</points>
<intersection>-79 12</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-79.5,-79,-79,-79</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<intersection>-79 9</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,-76.5,-51,-76.5</points>
<connection>
<GID>275</GID>
<name>IN_B_2</name></connection>
<intersection>-76.5 8</intersection>
<intersection>-70.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-70.5,-76.5,-70.5,-61.5</points>
<intersection>-76.5 1</intersection>
<intersection>-61.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-70.5,-61.5,-28.5,-61.5</points>
<connection>
<GID>273</GID>
<name>IN_B_2</name></connection>
<intersection>-70.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-76.5,-81,-76.5,-76.5</points>
<intersection>-81 9</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-79.5,-81,-76.5,-81</points>
<connection>
<GID>240</GID>
<name>OUT_2</name></connection>
<intersection>-76.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-77.5,-75.5,-51,-75.5</points>
<connection>
<GID>275</GID>
<name>IN_B_1</name></connection>
<intersection>-77.5 10</intersection>
<intersection>-71.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-71.5,-75.5,-71.5,-60.5</points>
<intersection>-75.5 1</intersection>
<intersection>-60.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-71.5,-60.5,-28.5,-60.5</points>
<connection>
<GID>273</GID>
<name>IN_B_1</name></connection>
<intersection>-71.5 8</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-77.5,-80,-77.5,-75.5</points>
<intersection>-80 14</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-79.5,-80,-77.5,-80</points>
<connection>
<GID>240</GID>
<name>OUT_1</name></connection>
<intersection>-77.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>347,-28,362.5,-28</points>
<connection>
<GID>241</GID>
<name>carry_out</name></connection>
<connection>
<GID>283</GID>
<name>carry_in</name></connection>
<intersection>348 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>348,-46.5,348,-28</points>
<connection>
<GID>400</GID>
<name>IN_1</name></connection>
<intersection>-28 1</intersection></vsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353.5,-67.5,353.5,-48</points>
<intersection>-67.5 1</intersection>
<intersection>-54.5 14</intersection>
<intersection>-48 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353.5,-67.5,370,-67.5</points>
<intersection>353.5 0</intersection>
<intersection>370 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>370,-73,370,-67.5</points>
<intersection>-73 3</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>368.5,-73,370,-73</points>
<connection>
<GID>302</GID>
<name>carry_in</name></connection>
<intersection>370 2</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>353.5,-48,364,-48</points>
<intersection>353.5 0</intersection>
<intersection>363 12</intersection>
<intersection>364 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>364,-49,364,-48</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<intersection>-48 8</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>363,-49,363,-48</points>
<connection>
<GID>288</GID>
<name>IN_2</name></connection>
<intersection>-48 8</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>349,-54.5,353.5,-54.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>349 18</intersection>
<intersection>353.5 0</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>349,-54.5,349,-52.5</points>
<connection>
<GID>400</GID>
<name>OUT</name></connection>
<intersection>-54.5 14</intersection></vsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>368,-69,368,-66.5</points>
<intersection>-69 3</intersection>
<intersection>-66.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>371.5,-66.5,371.5,-66</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>368,-66.5,371.5,-66.5</points>
<intersection>368 0</intersection>
<intersection>371.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>365.5,-69,368,-69</points>
<intersection>365.5 4</intersection>
<intersection>368 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>365.5,-70,365.5,-69</points>
<connection>
<GID>302</GID>
<name>IN_B_0</name></connection>
<intersection>-69 3</intersection></vsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>364.5,-70,364.5,-68.5</points>
<connection>
<GID>302</GID>
<name>IN_B_1</name></connection>
<intersection>-68.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>367.5,-68.5,367.5,-66</points>
<connection>
<GID>300</GID>
<name>OUT</name></connection>
<intersection>-68.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>364.5,-68.5,367.5,-68.5</points>
<intersection>364.5 0</intersection>
<intersection>367.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363.5,-70,363.5,-66</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<connection>
<GID>302</GID>
<name>IN_B_2</name></connection></vsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361,-69,361,-66</points>
<intersection>-69 3</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>359.5,-66,361,-66</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<intersection>361 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>361,-69,362.5,-69</points>
<intersection>361 0</intersection>
<intersection>362.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>362.5,-70,362.5,-69</points>
<connection>
<GID>302</GID>
<name>IN_B_3</name></connection>
<intersection>-69 3</intersection></vsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-74,-77.5,-51,-77.5</points>
<connection>
<GID>275</GID>
<name>IN_B_3</name></connection>
<intersection>-74 8</intersection>
<intersection>-69 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-69,-77.5,-69,-62.5</points>
<intersection>-77.5 1</intersection>
<intersection>-62.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-69,-62.5,-28.5,-62.5</points>
<connection>
<GID>273</GID>
<name>IN_B_3</name></connection>
<intersection>-69 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-74,-82,-74,-77.5</points>
<intersection>-82 9</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-79.5,-82,-74,-82</points>
<connection>
<GID>240</GID>
<name>OUT_3</name></connection>
<intersection>-74 8</intersection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>358.5,-60,358.5,-57</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>358.5,-57,365.5,-57</points>
<connection>
<GID>288</GID>
<name>OUT_3</name></connection>
<intersection>358.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,-57.5,366.5,-57</points>
<connection>
<GID>288</GID>
<name>OUT_2</name></connection>
<intersection>-57.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>362.5,-60,362.5,-57.5</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>362.5,-57.5,366.5,-57.5</points>
<intersection>362.5 1</intersection>
<intersection>366.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,-60,366.5,-58</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>367.5,-58,367.5,-57</points>
<connection>
<GID>288</GID>
<name>OUT_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>366.5,-58,367.5,-58</points>
<intersection>366.5 0</intersection>
<intersection>367.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370.5,-60,370.5,-58</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>368.5,-58,368.5,-57</points>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>368.5,-58,370.5,-58</points>
<intersection>368.5 1</intersection>
<intersection>370.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520.5,-4.5,520.5,-1</points>
<intersection>-4.5 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,-4.5,520.5,-4.5</points>
<connection>
<GID>325</GID>
<name>OUT_0</name></connection>
<intersection>520.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>520.5,-1,528,-1</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<intersection>520.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>513.5,8.5,528,8.5</points>
<connection>
<GID>406</GID>
<name>IN_1</name></connection>
<connection>
<GID>313</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>521,9.5,521,13</points>
<intersection>9.5 1</intersection>
<intersection>13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,9.5,521,9.5</points>
<connection>
<GID>313</GID>
<name>OUT_2</name></connection>
<intersection>521 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>521,13,528,13</points>
<connection>
<GID>405</GID>
<name>IN_1</name></connection>
<intersection>521 0</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>519.5,10.5,519.5,18.5</points>
<intersection>10.5 1</intersection>
<intersection>18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,10.5,519.5,10.5</points>
<connection>
<GID>313</GID>
<name>OUT_1</name></connection>
<intersection>519.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>519.5,18.5,528,18.5</points>
<connection>
<GID>404</GID>
<name>IN_1</name></connection>
<intersection>519.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520,11.5,520,29.5</points>
<intersection>11.5 1</intersection>
<intersection>29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,11.5,520,11.5</points>
<connection>
<GID>313</GID>
<name>OUT_0</name></connection>
<intersection>520 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>520,29.5,528,29.5</points>
<connection>
<GID>403</GID>
<name>IN_1</name></connection>
<intersection>520 0</intersection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509.5,20.5,509.5,22</points>
<connection>
<GID>312</GID>
<name>carry_out</name></connection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>509.5,20.5,528,20.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>509.5 0</intersection>
<intersection>525 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>525,-11,525,31.5</points>
<intersection>-11 33</intersection>
<intersection>-7 31</intersection>
<intersection>-3 30</intersection>
<intersection>1 29</intersection>
<intersection>10.5 3</intersection>
<intersection>15 6</intersection>
<intersection>20.5 1</intersection>
<intersection>31.5 28</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>525,10.5,528,10.5</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>525,15,528,15</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>525,31.5,528,31.5</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>525,1,528,1</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>525,-3,528,-3</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>525,-7,528,-7</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>525,-11,528,-11</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>525 2</intersection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>534,30.5,545.5,30.5</points>
<connection>
<GID>403</GID>
<name>OUT</name></connection>
<connection>
<GID>411</GID>
<name>IN_B_0</name></connection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51,-84.5,-51,-84.5</points>
<connection>
<GID>275</GID>
<name>IN_3</name></connection>
<connection>
<GID>285</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88,-52,-88,-44.5</points>
<intersection>-52 1</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-137,-52,-88,-52</points>
<intersection>-137 3</intersection>
<intersection>-88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-88,-44.5,-87.5,-44.5</points>
<connection>
<GID>236</GID>
<name>IN_2</name></connection>
<intersection>-88 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-137,-52,-137,-47.5</points>
<intersection>-52 1</intersection>
<intersection>-47.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-137.5,-47.5,-137,-47.5</points>
<connection>
<GID>232</GID>
<name>OUT_2</name></connection>
<intersection>-137 3</intersection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-137,-51,-87.5,-51</points>
<intersection>-137 3</intersection>
<intersection>-87.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-87.5,-51,-87.5,-45.5</points>
<connection>
<GID>236</GID>
<name>IN_3</name></connection>
<intersection>-51 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>-137,-51,-137,-45.5</points>
<intersection>-51 1</intersection>
<intersection>-45.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-137.5,-45.5,-137,-45.5</points>
<connection>
<GID>232</GID>
<name>OUT_3</name></connection>
<intersection>-137 3</intersection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-1,-77,-1,-77</points>
<connection>
<GID>304</GID>
<name>N_in2</name></connection>
<connection>
<GID>317</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-1,-79,-1,-79</points>
<connection>
<GID>317</GID>
<name>N_in2</name></connection>
<connection>
<GID>318</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>537.5,19.5,537.5,29.5</points>
<intersection>19.5 2</intersection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>537.5,29.5,545.5,29.5</points>
<connection>
<GID>411</GID>
<name>IN_B_1</name></connection>
<intersection>537.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>534,19.5,537.5,19.5</points>
<connection>
<GID>404</GID>
<name>OUT</name></connection>
<intersection>537.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84.5,-72.5,-84.5,-48.5</points>
<connection>
<GID>240</GID>
<name>carry_in</name></connection>
<connection>
<GID>236</GID>
<name>carry_out</name></connection>
<intersection>-55 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-84.5,-55,-75.5,-55</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<intersection>-84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-29,-5.5,-26</points>
<connection>
<GID>305</GID>
<name>IN_3</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-29,-5.5,-29</points>
<connection>
<GID>242</GID>
<name>OUT_3</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-28,-5.5,-27</points>
<connection>
<GID>305</GID>
<name>IN_2</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-28,-5.5,-28</points>
<connection>
<GID>242</GID>
<name>OUT_2</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-5.5,-28,-5.5,-27</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>-27 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-20.5,-27,-5.5,-27</points>
<connection>
<GID>242</GID>
<name>OUT_1</name></connection>
<intersection>-5.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-29,-5.5,-26</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-26,-5.5,-26</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-48.5,-52.5,-46,-52.5</points>
<intersection>-48.5 6</intersection>
<intersection>-46 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-48.5,-52.5,-48.5,-52</points>
<connection>
<GID>252</GID>
<name>A_less_B</name></connection>
<intersection>-52.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-46,-52.5,-46,-52</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>-52.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-66,-4,-63</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-63,-4,-63</points>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-65,-21,-64</points>
<intersection>-65 1</intersection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-65,-4,-65</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-64,-20.5,-64</points>
<connection>
<GID>273</GID>
<name>OUT_1</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-65,-4,-64</points>
<connection>
<GID>309</GID>
<name>IN_2</name></connection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-65,-4,-65</points>
<connection>
<GID>273</GID>
<name>OUT_2</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-66,-3.5,-63</points>
<intersection>-66 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-66,-3.5,-66</points>
<connection>
<GID>273</GID>
<name>OUT_3</name></connection>
<intersection>-3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-63,-3.5,-63</points>
<connection>
<GID>309</GID>
<name>IN_3</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45,-90,-45,-87.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<connection>
<GID>275</GID>
<name>A_less_B</name></connection></vsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-81,-1,-81</points>
<connection>
<GID>319</GID>
<name>N_in3</name></connection>
<connection>
<GID>318</GID>
<name>N_in2</name></connection>
<intersection>-1.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1.5,-81,-1.5,-80</points>
<intersection>-81 1</intersection>
<intersection>-80 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-2,-80,-1.5,-80</points>
<connection>
<GID>318</GID>
<name>N_in0</name></connection>
<intersection>-1.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,-56.5,-25.5,-35.5</points>
<connection>
<GID>273</GID>
<name>carry_in</name></connection>
<connection>
<GID>242</GID>
<name>carry_out</name></connection>
<intersection>-55.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-63.5,-55.5,-25.5,-55.5</points>
<intersection>-63.5 9</intersection>
<intersection>-25.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-63.5,-82.5,-63.5,-55.5</points>
<intersection>-82.5 10</intersection>
<intersection>-55.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-63.5,-82.5,-58.5,-82.5</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>-63.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-58.5,-80.5,-58.5,-80.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>316</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-52.5,-81.5,-51,-81.5</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<connection>
<GID>275</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-75,4.5,-11</points>
<intersection>-75 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-82.5,-11,4.5,-11</points>
<connection>
<GID>320</GID>
<name>OUT</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,-75,4.5,-75</points>
<connection>
<GID>304</GID>
<name>N_in3</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45,-46,-45,-33.5</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>-37.5 21</intersection>
<intersection>-33.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-45,-33.5,-36,-33.5</points>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<intersection>-45 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-45,-37.5,-36,-37.5</points>
<connection>
<GID>323</GID>
<name>IN_1</name></connection>
<intersection>-45 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-36.5,-29,-31.5</points>
<intersection>-36.5 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,-31.5,-28.5,-31.5</points>
<connection>
<GID>242</GID>
<name>IN_2</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-30,-36.5,-29,-36.5</points>
<connection>
<GID>323</GID>
<name>OUT</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-32.5,-29.5,-30.5</points>
<intersection>-32.5 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-30.5,-28.5,-30.5</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-30,-32.5,-29.5,-32.5</points>
<connection>
<GID>322</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-29.5,-29.5,-28.5</points>
<intersection>-29.5 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-29.5,-28.5,-29.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-30,-28.5,-29.5,-28.5</points>
<connection>
<GID>321</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-40.5,-28.5,-32.5</points>
<connection>
<GID>242</GID>
<name>IN_3</name></connection>
<intersection>-40.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-30,-40.5,-28.5,-40.5</points>
<connection>
<GID>324</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>538.5,14,538.5,28.5</points>
<intersection>14 1</intersection>
<intersection>28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534,14,538.5,14</points>
<connection>
<GID>405</GID>
<name>OUT</name></connection>
<intersection>538.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>538.5,28.5,545.5,28.5</points>
<connection>
<GID>411</GID>
<name>IN_B_2</name></connection>
<intersection>538.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-29.5,-36,-29.5</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<connection>
<GID>321</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-41.5,-36,-41.5</points>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<connection>
<GID>324</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-81.5,-38,-69.5</points>
<intersection>-81.5 28</intersection>
<intersection>-73.5 21</intersection>
<intersection>-69.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-38,-69.5,-35.5,-69.5</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>-38 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-38,-73.5,-35.5,-73.5</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<intersection>-38 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-38,-81.5,-36,-81.5</points>
<connection>
<GID>329</GID>
<name>OUT</name></connection>
<intersection>-38 0</intersection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-65.5,-35.5,-65.5</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<connection>
<GID>229</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-77.5,-35.5,-77.5</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<connection>
<GID>234</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539.5,9.5,539.5,27.5</points>
<intersection>9.5 2</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>539.5,27.5,545.5,27.5</points>
<connection>
<GID>411</GID>
<name>IN_B_3</name></connection>
<intersection>539.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>534,9.5,539.5,9.5</points>
<connection>
<GID>406</GID>
<name>OUT</name></connection>
<intersection>539.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-105.5,-77.5,-105.5,-16.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<connection>
<GID>271</GID>
<name>OUT</name></connection>
<intersection>-36.5 101</intersection>
<intersection>-32.5 39</intersection>
<intersection>-28.5 29</intersection>
<intersection>-24.5 28</intersection>
<intersection>-16.5 30</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-105.5,-24.5,-104.5,-24.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-105.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-105.5,-28.5,-104.5,-28.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-105.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-105.5,-16.5,-25.5,-16.5</points>
<intersection>-105.5 0</intersection>
<intersection>-84.5 233</intersection>
<intersection>-40 37</intersection>
<intersection>-25.5 226</intersection></hsegment>
<vsegment>
<ID>37</ID>
<points>-40,-88,-40,-16.5</points>
<intersection>-88 240</intersection>
<intersection>-75.5 90</intersection>
<intersection>-71.5 98</intersection>
<intersection>-67.5 95</intersection>
<intersection>-63.5 96</intersection>
<intersection>-39.5 237</intersection>
<intersection>-35.5 48</intersection>
<intersection>-31.5 45</intersection>
<intersection>-27.5 228</intersection>
<intersection>-16.5 30</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>-105.5,-32.5,-104.5,-32.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>-105.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>-40,-31.5,-36,-31.5</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-40,-35.5,-36,-35.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>90</ID>
<points>-40,-75.5,-35.5,-75.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>95</ID>
<points>-40,-67.5,-35.5,-67.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>96</ID>
<points>-40,-63.5,-35.5,-63.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>98</ID>
<points>-40,-71.5,-35.5,-71.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>101</ID>
<points>-105.5,-36.5,-104.5,-36.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>-105.5 0</intersection></hsegment>
<vsegment>
<ID>226</ID>
<points>-25.5,-19.5,-25.5,-16.5</points>
<connection>
<GID>242</GID>
<name>carry_in</name></connection>
<intersection>-16.5 30</intersection></vsegment>
<hsegment>
<ID>228</ID>
<points>-40,-27.5,-36,-27.5</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<vsegment>
<ID>233</ID>
<points>-84.5,-53,-84.5,-16.5</points>
<connection>
<GID>236</GID>
<name>carry_in</name></connection>
<intersection>-53 234</intersection>
<intersection>-16.5 30</intersection></vsegment>
<hsegment>
<ID>234</ID>
<points>-84.5,-53,-75.5,-53</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>-84.5 233</intersection></hsegment>
<hsegment>
<ID>237</ID>
<points>-40,-39.5,-36,-39.5</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>-40 37</intersection></hsegment>
<hsegment>
<ID>240</ID>
<points>-40,-88,-37,-88</points>
<intersection>-40 37</intersection>
<intersection>-37 241</intersection></hsegment>
<vsegment>
<ID>241</ID>
<points>-37,-88,-37,-87.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>-88 240</intersection></vsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>537,0,537,8.5</points>
<intersection>0 1</intersection>
<intersection>8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534,0,537,0</points>
<connection>
<GID>407</GID>
<name>OUT</name></connection>
<intersection>537 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>537,8.5,545.5,8.5</points>
<connection>
<GID>412</GID>
<name>IN_B_0</name></connection>
<intersection>537 0</intersection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>536,-4,536,7.5</points>
<intersection>-4 1</intersection>
<intersection>7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534,-4,536,-4</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>536 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>536,7.5,545.5,7.5</points>
<connection>
<GID>412</GID>
<name>IN_B_1</name></connection>
<intersection>536 0</intersection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>538,-8,538,6.5</points>
<intersection>-8 1</intersection>
<intersection>6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534,-8,538,-8</points>
<connection>
<GID>409</GID>
<name>OUT</name></connection>
<intersection>538 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>538,6.5,545.5,6.5</points>
<connection>
<GID>412</GID>
<name>IN_B_2</name></connection>
<intersection>538 0</intersection></hsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-76.5,-28.5,-69.5</points>
<connection>
<GID>273</GID>
<name>IN_3</name></connection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,-76.5,-28.5,-76.5</points>
<connection>
<GID>234</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539.5,-12,539.5,5.5</points>
<intersection>-12 3</intersection>
<intersection>5.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>534,-12,539.5,-12</points>
<connection>
<GID>410</GID>
<name>OUT</name></connection>
<intersection>539.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>539.5,5.5,545.5,5.5</points>
<connection>
<GID>412</GID>
<name>IN_B_3</name></connection>
<intersection>539.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-66.5,-29,-64.5</points>
<intersection>-66.5 1</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,-66.5,-28.5,-66.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,-64.5,-29,-64.5</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-68.5,-29.5,-67.5</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-67.5,-28.5,-67.5</points>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>538,-14.5,545.5,-14.5</points>
<intersection>538 3</intersection>
<intersection>545.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>538,-18,538,-14.5</points>
<connection>
<GID>311</GID>
<name>OUT_7</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>545.5,-14.5,545.5,-1.5</points>
<connection>
<GID>412</GID>
<name>IN_3</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-38.5,-106.5,-32</points>
<intersection>-38.5 5</intersection>
<intersection>-32 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-110.5,-32,-106.5,-32</points>
<connection>
<GID>227</GID>
<name>OUT_3</name></connection>
<intersection>-106.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106.5,-38.5,-104.5,-38.5</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-34.5,-106.5,-34</points>
<intersection>-34.5 5</intersection>
<intersection>-34 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-110.5,-34,-106.5,-34</points>
<connection>
<GID>227</GID>
<name>OUT_2</name></connection>
<intersection>-106.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106.5,-34.5,-104.5,-34.5</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-36,-106.5,-30.5</points>
<intersection>-36 4</intersection>
<intersection>-30.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-110.5,-36,-106.5,-36</points>
<connection>
<GID>227</GID>
<name>OUT_1</name></connection>
<intersection>-106.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106.5,-30.5,-104.5,-30.5</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-38,-106.5,-26.5</points>
<intersection>-38 4</intersection>
<intersection>-26.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-110.5,-38,-106.5,-38</points>
<connection>
<GID>227</GID>
<name>OUT_0</name></connection>
<intersection>-106.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106.5,-26.5,-104.5,-26.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>541.5,-19,541.5,-0.5</points>
<intersection>-19 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-19,541.5,-19</points>
<connection>
<GID>311</GID>
<name>OUT_6</name></connection>
<intersection>541.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>541.5,-0.5,545.5,-0.5</points>
<connection>
<GID>412</GID>
<name>IN_2</name></connection>
<intersection>541.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>542,-20,542,0.5</points>
<intersection>-20 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-20,542,-20</points>
<connection>
<GID>311</GID>
<name>OUT_5</name></connection>
<intersection>542 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>542,0.5,545.5,0.5</points>
<connection>
<GID>412</GID>
<name>IN_1</name></connection>
<intersection>542 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-21,540.5,1.5</points>
<intersection>-21 1</intersection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-21,540.5,-21</points>
<connection>
<GID>311</GID>
<name>OUT_4</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,1.5,545.5,1.5</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>540.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>544.5,-22,544.5,20.5</points>
<intersection>-22 1</intersection>
<intersection>20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-22,544.5,-22</points>
<connection>
<GID>311</GID>
<name>OUT_3</name></connection>
<intersection>544.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>544.5,20.5,545.5,20.5</points>
<connection>
<GID>411</GID>
<name>IN_3</name></connection>
<intersection>544.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107.5,-79.5,-107.5,-73</points>
<intersection>-79.5 3</intersection>
<intersection>-73 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-107.5,-79.5,-105.5,-79.5</points>
<connection>
<GID>226</GID>
<name>IN_1</name></connection>
<intersection>-107.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-112,-73,-107.5,-73</points>
<connection>
<GID>235</GID>
<name>OUT_3</name></connection>
<intersection>-107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107.5,-75.5,-107.5,-75</points>
<intersection>-75.5 3</intersection>
<intersection>-75 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-107.5,-75.5,-105.5,-75.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>-107.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-112,-75,-107.5,-75</points>
<connection>
<GID>235</GID>
<name>OUT_2</name></connection>
<intersection>-107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107.5,-77,-107.5,-71.5</points>
<intersection>-77 4</intersection>
<intersection>-71.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-107.5,-71.5,-105.5,-71.5</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>-107.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-112,-77,-107.5,-77</points>
<connection>
<GID>235</GID>
<name>OUT_1</name></connection>
<intersection>-107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107.5,-79,-107.5,-67.5</points>
<intersection>-79 4</intersection>
<intersection>-67.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-107.5,-67.5,-105.5,-67.5</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>-107.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-112,-79,-107.5,-79</points>
<connection>
<GID>235</GID>
<name>OUT_0</name></connection>
<intersection>-107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84.5,-92,-84.5,-88.5</points>
<connection>
<GID>240</GID>
<name>carry_out</name></connection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-84.5,-92,-45,-92</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>-84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93,-35.5,-93,-25.5</points>
<intersection>-35.5 1</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93,-35.5,-87.5,-35.5</points>
<connection>
<GID>236</GID>
<name>IN_B_0</name></connection>
<intersection>-93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-98.5,-25.5,-93,-25.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>-93 0</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93,-36.5,-93,-29.5</points>
<intersection>-36.5 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-98.5,-29.5,-93,-29.5</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>-93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-93,-36.5,-87.5,-36.5</points>
<connection>
<GID>236</GID>
<name>IN_B_1</name></connection>
<intersection>-93 0</intersection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93,-37.5,-93,-33.5</points>
<intersection>-37.5 1</intersection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93,-37.5,-87.5,-37.5</points>
<connection>
<GID>236</GID>
<name>IN_B_2</name></connection>
<intersection>-93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-98.5,-33.5,-93,-33.5</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>-93 0</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93,-38.5,-93,-37.5</points>
<intersection>-38.5 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-98.5,-37.5,-93,-37.5</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>-93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-93,-38.5,-87.5,-38.5</points>
<connection>
<GID>236</GID>
<name>IN_B_3</name></connection>
<intersection>-93 0</intersection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93.5,-75.5,-93.5,-66.5</points>
<intersection>-75.5 1</intersection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93.5,-75.5,-87.5,-75.5</points>
<connection>
<GID>240</GID>
<name>IN_B_0</name></connection>
<intersection>-93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-99.5,-66.5,-93.5,-66.5</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>-93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93.5,-76.5,-93.5,-70.5</points>
<intersection>-76.5 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-99.5,-70.5,-93.5,-70.5</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<intersection>-93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-93.5,-76.5,-87.5,-76.5</points>
<connection>
<GID>240</GID>
<name>IN_B_1</name></connection>
<intersection>-93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93.5,-77.5,-93.5,-74.5</points>
<intersection>-77.5 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93.5,-77.5,-87.5,-77.5</points>
<connection>
<GID>240</GID>
<name>IN_B_2</name></connection>
<intersection>-93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-99.5,-74.5,-93.5,-74.5</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<intersection>-93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-99.5,-78.5,-87.5,-78.5</points>
<connection>
<GID>226</GID>
<name>OUT</name></connection>
<connection>
<GID>240</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-54,-44,-52</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,-54,-44,-54</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>543.5,-23,543.5,21.5</points>
<intersection>-23 1</intersection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-23,543.5,-23</points>
<connection>
<GID>311</GID>
<name>OUT_2</name></connection>
<intersection>543.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>543.5,21.5,545.5,21.5</points>
<connection>
<GID>411</GID>
<name>IN_2</name></connection>
<intersection>543.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>542.5,-24,542.5,22.5</points>
<intersection>-24 1</intersection>
<intersection>22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-24,542.5,-24</points>
<connection>
<GID>311</GID>
<name>OUT_1</name></connection>
<intersection>542.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>542.5,22.5,545.5,22.5</points>
<connection>
<GID>411</GID>
<name>IN_1</name></connection>
<intersection>542.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>541,-25,541,23.5</points>
<intersection>-25 1</intersection>
<intersection>23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>538,-25,541,-25</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<intersection>541 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>541,23.5,545.5,23.5</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>541 0</intersection></hsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-91,-35,-87.5</points>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-91,-35,-91</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,-12.5,-268,-12</points>
<connection>
<GID>356</GID>
<name>IN_1</name></connection>
<connection>
<GID>354</GID>
<name>OUT_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-268,-12,-250,-12</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-266,-14,-266,-12.5</points>
<connection>
<GID>337</GID>
<name>OUT_0</name></connection>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-266,-14,-250,-14</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<intersection>-266 0</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-241,-41,-216,-41</points>
<connection>
<GID>343</GID>
<name>OUT_0</name></connection>
<connection>
<GID>350</GID>
<name>IN_B_0</name></connection>
<intersection>-236.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-236.5,-41,-236.5,-24.5</points>
<intersection>-41 1</intersection>
<intersection>-24.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-236.5,-24.5,-190,-24.5</points>
<connection>
<GID>346</GID>
<name>IN_B_0</name></connection>
<intersection>-236.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-241,-43,-216,-43</points>
<connection>
<GID>343</GID>
<name>OUT_2</name></connection>
<connection>
<GID>350</GID>
<name>IN_B_2</name></connection>
<intersection>-234.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-234.5,-43,-234.5,-26.5</points>
<intersection>-43 1</intersection>
<intersection>-26.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-234.5,-26.5,-190,-26.5</points>
<connection>
<GID>346</GID>
<name>IN_B_2</name></connection>
<intersection>-234.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-241,-42,-216,-42</points>
<connection>
<GID>343</GID>
<name>OUT_1</name></connection>
<connection>
<GID>350</GID>
<name>IN_B_1</name></connection>
<intersection>-235.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-235.5,-42,-235.5,-25.5</points>
<intersection>-42 1</intersection>
<intersection>-25.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-235.5,-25.5,-190,-25.5</points>
<connection>
<GID>346</GID>
<name>IN_B_1</name></connection>
<intersection>-235.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-241,-44,-216,-44</points>
<connection>
<GID>343</GID>
<name>OUT_3</name></connection>
<connection>
<GID>350</GID>
<name>IN_B_3</name></connection>
<intersection>-233 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-233,-44,-233,-27.5</points>
<intersection>-44 1</intersection>
<intersection>-27.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-233,-27.5,-190,-27.5</points>
<connection>
<GID>346</GID>
<name>IN_B_3</name></connection>
<intersection>-233 6</intersection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-221,-51,-216,-51</points>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection>
<connection>
<GID>350</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-220.5,-48,-216,-48</points>
<connection>
<GID>352</GID>
<name>OUT_0</name></connection>
<connection>
<GID>350</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-298,-96,-249,-96</points>
<intersection>-298 5</intersection>
<intersection>-249 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-298,-96,-298,-88.5</points>
<connection>
<GID>344</GID>
<name>OUT_3</name></connection>
<intersection>-96 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-249,-96,-249,-87.5</points>
<connection>
<GID>345</GID>
<name>IN_3</name></connection>
<intersection>-96 1</intersection></vsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249,-96,-249,-86.5</points>
<connection>
<GID>345</GID>
<name>IN_2</name></connection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-298,-96,-249,-96</points>
<intersection>-298 3</intersection>
<intersection>-249 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-298,-96,-298,-90.5</points>
<connection>
<GID>344</GID>
<name>OUT_2</name></connection>
<intersection>-96 1</intersection></vsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249,-96,-249,-85.5</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-298,-96,-249,-96</points>
<intersection>-298 3</intersection>
<intersection>-249 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-298,-96,-298,-92.5</points>
<connection>
<GID>344</GID>
<name>OUT_1</name></connection>
<intersection>-96 1</intersection></vsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249,-96,-249,-84.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-298,-96,-249,-96</points>
<intersection>-298 3</intersection>
<intersection>-249 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-298,-96,-298,-94.5</points>
<connection>
<GID>344</GID>
<name>OUT_0</name></connection>
<intersection>-96 1</intersection></vsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249,-56.5,-249,-44.5</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-298.5,-56.5,-249,-56.5</points>
<intersection>-298.5 3</intersection>
<intersection>-249 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-298.5,-57,-298.5,-56.5</points>
<connection>
<GID>339</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249,-55,-249,-45.5</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<intersection>-55 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-298.5,-55,-249,-55</points>
<connection>
<GID>339</GID>
<name>OUT_1</name></connection>
<intersection>-249 0</intersection></hsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-240.5,-76.5,-214,-76.5</points>
<connection>
<GID>359</GID>
<name>IN_B_0</name></connection>
<intersection>-240.5 9</intersection>
<intersection>-234 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-234,-76.5,-234,-61.5</points>
<intersection>-76.5 1</intersection>
<intersection>-61.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-234,-61.5,-190,-61.5</points>
<connection>
<GID>358</GID>
<name>IN_B_0</name></connection>
<intersection>-234 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-240.5,-81,-240.5,-76.5</points>
<intersection>-81 12</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-241,-81,-240.5,-81</points>
<connection>
<GID>345</GID>
<name>OUT_0</name></connection>
<intersection>-240.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-238,-78.5,-214,-78.5</points>
<connection>
<GID>359</GID>
<name>IN_B_2</name></connection>
<intersection>-238 8</intersection>
<intersection>-232 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-232,-78.5,-232,-63.5</points>
<intersection>-78.5 1</intersection>
<intersection>-63.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-232,-63.5,-190,-63.5</points>
<connection>
<GID>358</GID>
<name>IN_B_2</name></connection>
<intersection>-232 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-238,-83,-238,-78.5</points>
<intersection>-83 9</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-241,-83,-238,-83</points>
<connection>
<GID>345</GID>
<name>OUT_2</name></connection>
<intersection>-238 8</intersection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-239,-77.5,-214,-77.5</points>
<connection>
<GID>359</GID>
<name>IN_B_1</name></connection>
<intersection>-239 10</intersection>
<intersection>-233 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-233,-77.5,-233,-62.5</points>
<intersection>-77.5 1</intersection>
<intersection>-62.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-233,-62.5,-190,-62.5</points>
<connection>
<GID>358</GID>
<name>IN_B_1</name></connection>
<intersection>-233 8</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-239,-82,-239,-77.5</points>
<intersection>-82 14</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-241,-82,-239,-82</points>
<connection>
<GID>345</GID>
<name>OUT_1</name></connection>
<intersection>-239 10</intersection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-235.5,-79.5,-214,-79.5</points>
<connection>
<GID>359</GID>
<name>IN_B_3</name></connection>
<intersection>-235.5 8</intersection>
<intersection>-230.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-230.5,-79.5,-230.5,-64.5</points>
<intersection>-79.5 1</intersection>
<intersection>-64.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-230.5,-64.5,-190,-64.5</points>
<connection>
<GID>358</GID>
<name>IN_B_3</name></connection>
<intersection>-230.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-235.5,-84,-235.5,-79.5</points>
<intersection>-84 9</intersection>
<intersection>-79.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-241,-84,-235.5,-84</points>
<connection>
<GID>345</GID>
<name>OUT_3</name></connection>
<intersection>-235.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-214.5,-86.5,-214,-86.5</points>
<connection>
<GID>361</GID>
<name>OUT_0</name></connection>
<connection>
<GID>359</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249.5,-50.5,-249.5,-46.5</points>
<intersection>-50.5 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-298.5,-50.5,-249.5,-50.5</points>
<intersection>-298.5 3</intersection>
<intersection>-249.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-249.5,-46.5,-249,-46.5</points>
<connection>
<GID>343</GID>
<name>IN_2</name></connection>
<intersection>-249.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-298.5,-53,-298.5,-50.5</points>
<connection>
<GID>339</GID>
<name>OUT_2</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-298.5,-53,-249,-53</points>
<intersection>-298.5 3</intersection>
<intersection>-249 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-249,-53,-249,-47.5</points>
<connection>
<GID>343</GID>
<name>IN_3</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>-298.5,-53,-298.5,-51</points>
<connection>
<GID>339</GID>
<name>OUT_3</name></connection>
<intersection>-53 1</intersection></vsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-162.5,-79,-162.5,-79</points>
<connection>
<GID>362</GID>
<name>N_in2</name></connection>
<connection>
<GID>369</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-162.5,-81,-162.5,-81</points>
<connection>
<GID>369</GID>
<name>N_in2</name></connection>
<connection>
<GID>370</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-246,-67,-246,-50.5</points>
<connection>
<GID>343</GID>
<name>carry_out</name></connection>
<connection>
<GID>386</GID>
<name>IN_1</name></connection>
<intersection>-57 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-246,-57,-237,-57</points>
<connection>
<GID>377</GID>
<name>IN_1</name></connection>
<intersection>-246 0</intersection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-167,-31,-167,-28</points>
<connection>
<GID>363</GID>
<name>IN_3</name></connection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-31,-167,-31</points>
<connection>
<GID>346</GID>
<name>OUT_3</name></connection>
<intersection>-167 0</intersection></hsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-167,-30,-167,-29</points>
<connection>
<GID>363</GID>
<name>IN_2</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-30,-167,-30</points>
<connection>
<GID>346</GID>
<name>OUT_2</name></connection>
<intersection>-167 0</intersection></hsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-167,-30,-167,-29</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<intersection>-29 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-182,-29,-167,-29</points>
<connection>
<GID>346</GID>
<name>OUT_1</name></connection>
<intersection>-167 3</intersection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-167,-31,-167,-28</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-28,-167,-28</points>
<connection>
<GID>346</GID>
<name>OUT_0</name></connection>
<intersection>-167 0</intersection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-210,-54.5,-207.5,-54.5</points>
<intersection>-210 6</intersection>
<intersection>-207.5 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-210,-54.5,-210,-54</points>
<connection>
<GID>350</GID>
<name>A_less_B</name></connection>
<intersection>-54.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-207.5,-54.5,-207.5,-54</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-54.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-165.5,-68,-165.5,-65</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-65,-165.5,-65</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>-165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-182.5,-67,-182.5,-66</points>
<intersection>-67 1</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182.5,-67,-165.5,-67</points>
<connection>
<GID>365</GID>
<name>IN_1</name></connection>
<intersection>-182.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-182.5,-66,-182,-66</points>
<connection>
<GID>358</GID>
<name>OUT_1</name></connection>
<intersection>-182.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-165.5,-67,-165.5,-66</points>
<connection>
<GID>365</GID>
<name>IN_2</name></connection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-67,-165.5,-67</points>
<connection>
<GID>358</GID>
<name>OUT_2</name></connection>
<intersection>-165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-165,-68,-165,-65</points>
<intersection>-68 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-68,-165,-68</points>
<connection>
<GID>358</GID>
<name>OUT_3</name></connection>
<intersection>-165 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-165.5,-65,-165,-65</points>
<connection>
<GID>365</GID>
<name>IN_3</name></connection>
<intersection>-165 0</intersection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>533,-16,533,-15</points>
<connection>
<GID>311</GID>
<name>load</name></connection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>533.5,-15,533.5,-14.5</points>
<connection>
<GID>413</GID>
<name>OUT_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>533,-15,533.5,-15</points>
<intersection>533 0</intersection>
<intersection>533.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-163,-83,-162.5,-83</points>
<connection>
<GID>371</GID>
<name>N_in3</name></connection>
<connection>
<GID>370</GID>
<name>N_in2</name></connection>
<intersection>-163 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-163,-83,-163,-82</points>
<intersection>-83 1</intersection>
<intersection>-82 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-163.5,-82,-163,-82</points>
<connection>
<GID>370</GID>
<name>N_in0</name></connection>
<intersection>-163 4</intersection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-187,-58.5,-187,-37.5</points>
<connection>
<GID>346</GID>
<name>carry_out</name></connection>
<connection>
<GID>358</GID>
<name>carry_in</name></connection>
<intersection>-58.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-225,-58.5,-187,-58.5</points>
<intersection>-225 9</intersection>
<intersection>-187 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-225,-84.5,-225,-58.5</points>
<intersection>-84.5 10</intersection>
<intersection>-58.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-225,-84.5,-220,-84.5</points>
<connection>
<GID>367</GID>
<name>IN_1</name></connection>
<intersection>-225 9</intersection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-220,-82.5,-220,-82.5</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>567,-33.5,567,2</points>
<intersection>-33.5 5</intersection>
<intersection>2 13</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>524.5,-33.5,584,-33.5</points>
<connection>
<GID>310</GID>
<name>IN_7</name></connection>
<intersection>524.5 8</intersection>
<intersection>567 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>524.5,-33.5,524.5,-17</points>
<intersection>-33.5 5</intersection>
<intersection>-17 14</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>553.5,2,567,2</points>
<connection>
<GID>412</GID>
<name>OUT_3</name></connection>
<intersection>567 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>524.5,-17,530,-17</points>
<intersection>524.5 8</intersection>
<intersection>530 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>530,-18,530,-17</points>
<connection>
<GID>311</GID>
<name>IN_7</name></connection>
<intersection>-17 14</intersection></vsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-157,-77,-157,-13</points>
<intersection>-77 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-244,-13,-157,-13</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<intersection>-157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-162.5,-77,-157,-77</points>
<connection>
<GID>362</GID>
<name>N_in3</name></connection>
<intersection>-157 0</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-206.5,-48,-206.5,-35.5</points>
<connection>
<GID>364</GID>
<name>OUT</name></connection>
<intersection>-39.5 21</intersection>
<intersection>-35.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-206.5,-35.5,-197.5,-35.5</points>
<connection>
<GID>374</GID>
<name>IN_1</name></connection>
<intersection>-206.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-206.5,-39.5,-197.5,-39.5</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<intersection>-206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-190.5,-38.5,-190.5,-33.5</points>
<intersection>-38.5 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-190.5,-33.5,-190,-33.5</points>
<connection>
<GID>346</GID>
<name>IN_2</name></connection>
<intersection>-190.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-191.5,-38.5,-190.5,-38.5</points>
<connection>
<GID>375</GID>
<name>OUT</name></connection>
<intersection>-190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-191,-34.5,-191,-32.5</points>
<intersection>-34.5 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-191,-32.5,-190,-32.5</points>
<connection>
<GID>346</GID>
<name>IN_1</name></connection>
<intersection>-191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-191.5,-34.5,-191,-34.5</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<intersection>-191 0</intersection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-191,-31.5,-191,-30.5</points>
<intersection>-31.5 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-191,-31.5,-190,-31.5</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>-191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-191.5,-30.5,-191,-30.5</points>
<connection>
<GID>373</GID>
<name>OUT</name></connection>
<intersection>-191 0</intersection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-190,-42.5,-190,-34.5</points>
<connection>
<GID>346</GID>
<name>IN_3</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-191.5,-42.5,-190,-42.5</points>
<connection>
<GID>376</GID>
<name>OUT</name></connection>
<intersection>-190 0</intersection></hsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-197.5,-31.5,-197.5,-31.5</points>
<connection>
<GID>373</GID>
<name>IN_1</name></connection>
<connection>
<GID>379</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-197.5,-43.5,-197.5,-43.5</points>
<connection>
<GID>376</GID>
<name>IN_1</name></connection>
<connection>
<GID>380</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-199.5,-89.5,-199.5,-71.5</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>-75.5 21</intersection>
<intersection>-71.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-199.5,-71.5,-197,-71.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>-199.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-199.5,-75.5,-197,-75.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>-199.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-197,-67.5,-197,-67.5</points>
<connection>
<GID>336</GID>
<name>IN_1</name></connection>
<connection>
<GID>381</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-197,-79.5,-197,-79.5</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<connection>
<GID>341</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-270.5,-79.5,-270.5,-18.5</points>
<intersection>-79.5 246</intersection>
<intersection>-75.5 247</intersection>
<intersection>-71.5 248</intersection>
<intersection>-67.5 249</intersection>
<intersection>-38.5 101</intersection>
<intersection>-34.5 39</intersection>
<intersection>-30.5 29</intersection>
<intersection>-26.5 28</intersection>
<intersection>-18.5 30</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-270.5,-26.5,-266,-26.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-270.5,-30.5,-266,-30.5</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-270.5,-18.5,-187,-18.5</points>
<connection>
<GID>356</GID>
<name>OUT</name></connection>
<intersection>-270.5 0</intersection>
<intersection>-244 233</intersection>
<intersection>-202 37</intersection>
<intersection>-187 226</intersection></hsegment>
<vsegment>
<ID>37</ID>
<points>-202,-95.5,-202,-18.5</points>
<intersection>-95.5 255</intersection>
<intersection>-77.5 90</intersection>
<intersection>-73.5 98</intersection>
<intersection>-69.5 95</intersection>
<intersection>-65.5 96</intersection>
<intersection>-41.5 237</intersection>
<intersection>-37.5 48</intersection>
<intersection>-33.5 45</intersection>
<intersection>-29.5 228</intersection>
<intersection>-18.5 30</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>-270.5,-34.5,-266,-34.5</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>-202,-33.5,-197.5,-33.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-202,-37.5,-197.5,-37.5</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>90</ID>
<points>-202,-77.5,-197,-77.5</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>95</ID>
<points>-202,-69.5,-197,-69.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>96</ID>
<points>-202,-65.5,-197,-65.5</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>98</ID>
<points>-202,-73.5,-197,-73.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>101</ID>
<points>-270.5,-38.5,-266,-38.5</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<vsegment>
<ID>226</ID>
<points>-187,-21.5,-187,-18.5</points>
<connection>
<GID>346</GID>
<name>carry_in</name></connection>
<intersection>-18.5 30</intersection></vsegment>
<hsegment>
<ID>228</ID>
<points>-202,-29.5,-197.5,-29.5</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<vsegment>
<ID>233</ID>
<points>-244,-67,-244,-18.5</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>-55 234</intersection>
<intersection>-34.5 256</intersection>
<intersection>-18.5 30</intersection></vsegment>
<hsegment>
<ID>234</ID>
<points>-244,-55,-237,-55</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>-244 233</intersection></hsegment>
<hsegment>
<ID>237</ID>
<points>-202,-41.5,-197.5,-41.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>246</ID>
<points>-270.5,-79.5,-267,-79.5</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>247</ID>
<points>-270.5,-75.5,-267,-75.5</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>248</ID>
<points>-270.5,-71.5,-267,-71.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>249</ID>
<points>-270.5,-67.5,-267,-67.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>-270.5 0</intersection></hsegment>
<hsegment>
<ID>255</ID>
<points>-202,-95.5,-200.5,-95.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>-202 37</intersection></hsegment>
<hsegment>
<ID>256</ID>
<points>-246,-34.5,-244,-34.5</points>
<connection>
<GID>343</GID>
<name>carry_in</name></connection>
<intersection>-244 233</intersection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-190,-78.5,-190,-71.5</points>
<connection>
<GID>358</GID>
<name>IN_3</name></connection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-191,-78.5,-190,-78.5</points>
<connection>
<GID>341</GID>
<name>OUT</name></connection>
<intersection>-190 0</intersection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-190.5,-68.5,-190.5,-66.5</points>
<intersection>-68.5 1</intersection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-190.5,-68.5,-190,-68.5</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>-190.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-191,-66.5,-190.5,-66.5</points>
<connection>
<GID>336</GID>
<name>OUT</name></connection>
<intersection>-190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-191,-70.5,-191,-69.5</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-191,-69.5,-190,-69.5</points>
<connection>
<GID>358</GID>
<name>IN_1</name></connection>
<intersection>-191 0</intersection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-190.5,-74.5,-190.5,-70.5</points>
<intersection>-74.5 4</intersection>
<intersection>-70.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-190.5,-70.5,-190,-70.5</points>
<connection>
<GID>358</GID>
<name>IN_2</name></connection>
<intersection>-190.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-191,-74.5,-190.5,-74.5</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<intersection>-190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,-40.5,-268,-34</points>
<intersection>-40.5 5</intersection>
<intersection>-34 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-272,-34,-268,-34</points>
<connection>
<GID>335</GID>
<name>OUT_3</name></connection>
<intersection>-268 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-268,-40.5,-266,-40.5</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,-36.5,-268,-36</points>
<intersection>-36.5 5</intersection>
<intersection>-36 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-272,-36,-268,-36</points>
<connection>
<GID>335</GID>
<name>OUT_2</name></connection>
<intersection>-268 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-268,-36.5,-266,-36.5</points>
<connection>
<GID>357</GID>
<name>IN_1</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,-38,-268,-32.5</points>
<intersection>-38 4</intersection>
<intersection>-32.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-272,-38,-268,-38</points>
<connection>
<GID>335</GID>
<name>OUT_1</name></connection>
<intersection>-268 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-268,-32.5,-266,-32.5</points>
<connection>
<GID>348</GID>
<name>IN_1</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,-40,-268,-28.5</points>
<intersection>-40 4</intersection>
<intersection>-28.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-272,-40,-268,-40</points>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection>
<intersection>-268 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-268,-28.5,-266,-28.5</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-269,-81.5,-269,-75</points>
<intersection>-81.5 3</intersection>
<intersection>-75 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-269,-81.5,-267,-81.5</points>
<connection>
<GID>334</GID>
<name>IN_1</name></connection>
<intersection>-269 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-273.5,-75,-269,-75</points>
<connection>
<GID>342</GID>
<name>OUT_3</name></connection>
<intersection>-269 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-269,-77.5,-269,-77</points>
<intersection>-77.5 3</intersection>
<intersection>-77 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-269,-77.5,-267,-77.5</points>
<connection>
<GID>333</GID>
<name>IN_1</name></connection>
<intersection>-269 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-273.5,-77,-269,-77</points>
<connection>
<GID>342</GID>
<name>OUT_2</name></connection>
<intersection>-269 0</intersection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-269,-79,-269,-73.5</points>
<intersection>-79 4</intersection>
<intersection>-73.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-269,-73.5,-267,-73.5</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<intersection>-269 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-273.5,-79,-269,-79</points>
<connection>
<GID>342</GID>
<name>OUT_1</name></connection>
<intersection>-269 0</intersection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-269,-81,-269,-69.5</points>
<intersection>-81 4</intersection>
<intersection>-69.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-269,-69.5,-267,-69.5</points>
<connection>
<GID>331</GID>
<name>IN_1</name></connection>
<intersection>-269 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-273.5,-81,-269,-81</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<intersection>-269 0</intersection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-246,-98.5,-246,-90.5</points>
<connection>
<GID>345</GID>
<name>carry_out</name></connection>
<intersection>-98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-246,-98.5,-206.5,-98.5</points>
<connection>
<GID>366</GID>
<name>IN_1</name></connection>
<intersection>-246 0</intersection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-254.5,-37.5,-254.5,-27.5</points>
<intersection>-37.5 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-254.5,-37.5,-249,-37.5</points>
<connection>
<GID>343</GID>
<name>IN_B_0</name></connection>
<intersection>-254.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-260,-27.5,-254.5,-27.5</points>
<connection>
<GID>347</GID>
<name>OUT</name></connection>
<intersection>-254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-254.5,-38.5,-254.5,-31.5</points>
<intersection>-38.5 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-260,-31.5,-254.5,-31.5</points>
<connection>
<GID>348</GID>
<name>OUT</name></connection>
<intersection>-254.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-254.5,-38.5,-249,-38.5</points>
<connection>
<GID>343</GID>
<name>IN_B_1</name></connection>
<intersection>-254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-254.5,-39.5,-254.5,-35.5</points>
<intersection>-39.5 1</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-254.5,-39.5,-249,-39.5</points>
<connection>
<GID>343</GID>
<name>IN_B_2</name></connection>
<intersection>-254.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-260,-35.5,-254.5,-35.5</points>
<connection>
<GID>357</GID>
<name>OUT</name></connection>
<intersection>-254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-254.5,-40.5,-254.5,-39.5</points>
<intersection>-40.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-260,-39.5,-254.5,-39.5</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<intersection>-254.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-254.5,-40.5,-249,-40.5</points>
<connection>
<GID>343</GID>
<name>IN_B_3</name></connection>
<intersection>-254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-255,-77.5,-255,-68.5</points>
<intersection>-77.5 1</intersection>
<intersection>-68.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-255,-77.5,-249,-77.5</points>
<connection>
<GID>345</GID>
<name>IN_B_0</name></connection>
<intersection>-255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-261,-68.5,-255,-68.5</points>
<connection>
<GID>331</GID>
<name>OUT</name></connection>
<intersection>-255 0</intersection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-255,-78.5,-255,-72.5</points>
<intersection>-78.5 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-261,-72.5,-255,-72.5</points>
<connection>
<GID>332</GID>
<name>OUT</name></connection>
<intersection>-255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-255,-78.5,-249,-78.5</points>
<connection>
<GID>345</GID>
<name>IN_B_1</name></connection>
<intersection>-255 0</intersection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-255,-79.5,-255,-76.5</points>
<intersection>-79.5 1</intersection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-255,-79.5,-249,-79.5</points>
<connection>
<GID>345</GID>
<name>IN_B_2</name></connection>
<intersection>-255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-261,-76.5,-255,-76.5</points>
<connection>
<GID>333</GID>
<name>OUT</name></connection>
<intersection>-255 0</intersection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-261,-80.5,-249,-80.5</points>
<connection>
<GID>334</GID>
<name>OUT</name></connection>
<connection>
<GID>345</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-205.5,-56,-205.5,-54</points>
<connection>
<GID>364</GID>
<name>IN_1</name></connection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-231,-56,-205.5,-56</points>
<connection>
<GID>377</GID>
<name>OUT</name></connection>
<intersection>-205.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>564.5,-34.5,564.5,3</points>
<intersection>-34.5 1</intersection>
<intersection>3 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-34.5,584,-34.5</points>
<connection>
<GID>310</GID>
<name>IN_6</name></connection>
<intersection>527.5 6</intersection>
<intersection>564.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>527.5,-34.5,527.5,-19</points>
<intersection>-34.5 1</intersection>
<intersection>-19 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>553.5,3,564.5,3</points>
<connection>
<GID>412</GID>
<name>OUT_2</name></connection>
<intersection>564.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>527.5,-19,530,-19</points>
<connection>
<GID>311</GID>
<name>IN_6</name></connection>
<intersection>527.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-214,-83.5,-214,-83.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-198.5,-97.5,-198.5,-95.5</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-200.5,-97.5,-198.5,-97.5</points>
<connection>
<GID>366</GID>
<name>OUT</name></connection>
<intersection>-198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>561.5,-35.5,561.5,4</points>
<intersection>-35.5 1</intersection>
<intersection>4 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>526.5,-35.5,584,-35.5</points>
<connection>
<GID>310</GID>
<name>IN_5</name></connection>
<intersection>526.5 6</intersection>
<intersection>561.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>526.5,-35.5,526.5,-20</points>
<intersection>-35.5 1</intersection>
<intersection>-20 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>553.5,4,561.5,4</points>
<connection>
<GID>412</GID>
<name>OUT_1</name></connection>
<intersection>561.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>526.5,-20,530,-20</points>
<connection>
<GID>311</GID>
<name>IN_5</name></connection>
<intersection>526.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-172,-78,-172,-77.5</points>
<connection>
<GID>385</GID>
<name>N_in3</name></connection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-187,-78,-172,-78</points>
<intersection>-187 2</intersection>
<intersection>-172 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-187,-78,-187,-74.5</points>
<connection>
<GID>358</GID>
<name>carry_out</name></connection>
<intersection>-78 1</intersection></vsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>558.5,-36.5,558.5,5</points>
<intersection>-36.5 1</intersection>
<intersection>5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>529,-36.5,584,-36.5</points>
<connection>
<GID>310</GID>
<name>IN_4</name></connection>
<intersection>529 6</intersection>
<intersection>558.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>529,-36.5,529,-21</points>
<intersection>-36.5 1</intersection>
<intersection>-21 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>553.5,5,558.5,5</points>
<connection>
<GID>412</GID>
<name>OUT_0</name></connection>
<intersection>558.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>529,-21,530,-21</points>
<connection>
<GID>311</GID>
<name>IN_4</name></connection>
<intersection>529 6</intersection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>572.5,-37.5,572.5,24</points>
<intersection>-37.5 1</intersection>
<intersection>24 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>529.5,-37.5,584,-37.5</points>
<connection>
<GID>310</GID>
<name>IN_3</name></connection>
<intersection>529.5 6</intersection>
<intersection>572.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>529.5,-37.5,529.5,-22</points>
<intersection>-37.5 1</intersection>
<intersection>-22 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>553.5,24,572.5,24</points>
<connection>
<GID>411</GID>
<name>OUT_3</name></connection>
<intersection>572.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>529.5,-22,530,-22</points>
<connection>
<GID>311</GID>
<name>IN_3</name></connection>
<intersection>529.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-208,-96.5,-208,-89.5</points>
<connection>
<GID>359</GID>
<name>A_less_B</name></connection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-208,-96.5,-206.5,-96.5</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>-208 0</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-162.5,-84,-162.5,-80</points>
<intersection>-84 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-162.5,-84,-161.5,-84</points>
<connection>
<GID>371</GID>
<name>N_in1</name></connection>
<intersection>-162.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-163.5,-80,-162.5,-80</points>
<connection>
<GID>369</GID>
<name>N_in0</name></connection>
<intersection>-162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-245,-74.5,-245,-73</points>
<connection>
<GID>386</GID>
<name>OUT</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-246,-74.5,-245,-74.5</points>
<connection>
<GID>345</GID>
<name>carry_in</name></connection>
<intersection>-245 0</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-81.5,359,-78</points>
<connection>
<GID>302</GID>
<name>OUT_3</name></connection>
<intersection>-81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-81.5,364,-81.5</points>
<connection>
<GID>308</GID>
<name>IN_3</name></connection>
<intersection>359 0</intersection></hsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>360,-82.5,360,-78</points>
<connection>
<GID>302</GID>
<name>OUT_2</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360,-82.5,364,-82.5</points>
<connection>
<GID>308</GID>
<name>IN_2</name></connection>
<intersection>360 0</intersection></hsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361,-83.5,361,-78</points>
<connection>
<GID>302</GID>
<name>OUT_1</name></connection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361,-83.5,364,-83.5</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>361 0</intersection></hsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362,-84.5,362,-78</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>362,-84.5,364,-84.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>362 0</intersection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>314.5,-58.5,339,-58.5</points>
<intersection>314.5 26</intersection>
<intersection>327 39</intersection>
<intersection>331 27</intersection>
<intersection>335 28</intersection>
<intersection>339 29</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>314.5,-82.5,314.5,-56.5</points>
<connection>
<GID>397</GID>
<name>OUT_0</name></connection>
<intersection>-82.5 40</intersection>
<intersection>-69 30</intersection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>331,-60,331,-58.5</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>335,-60,335,-58.5</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>339,-60,339,-58.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>314.5,-69,324,-69</points>
<intersection>314.5 26</intersection>
<intersection>322 42</intersection>
<intersection>324 32</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>324,-70,324,-69</points>
<connection>
<GID>391</GID>
<name>IN_1</name></connection>
<intersection>-69 30</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>327,-60,327,-58.5</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>40</ID>
<points>314.5,-82.5,317,-82.5</points>
<connection>
<GID>396</GID>
<name>N_in0</name></connection>
<intersection>314.5 26</intersection></hsegment>
<vsegment>
<ID>42</ID>
<points>322,-70,322,-69</points>
<connection>
<GID>391</GID>
<name>IN_3</name></connection>
<intersection>-69 30</intersection></vsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334.5,-69,334.5,-66.5</points>
<intersection>-69 3</intersection>
<intersection>-66.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>338,-66.5,338,-66</points>
<connection>
<GID>390</GID>
<name>OUT</name></connection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>334.5,-66.5,338,-66.5</points>
<intersection>334.5 0</intersection>
<intersection>338 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>332,-69,334.5,-69</points>
<intersection>332 4</intersection>
<intersection>334.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>332,-70,332,-69</points>
<connection>
<GID>391</GID>
<name>IN_B_0</name></connection>
<intersection>-69 3</intersection></vsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331,-70,331,-68.5</points>
<connection>
<GID>391</GID>
<name>IN_B_1</name></connection>
<intersection>-68.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>334,-68.5,334,-66</points>
<connection>
<GID>389</GID>
<name>OUT</name></connection>
<intersection>-68.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>331,-68.5,334,-68.5</points>
<intersection>331 0</intersection>
<intersection>334 1</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,-70,330,-66</points>
<connection>
<GID>388</GID>
<name>OUT</name></connection>
<connection>
<GID>391</GID>
<name>IN_B_2</name></connection></vsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327.5,-69,327.5,-66</points>
<intersection>-69 3</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>326,-66,327.5,-66</points>
<connection>
<GID>387</GID>
<name>OUT</name></connection>
<intersection>327.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>327.5,-69,329,-69</points>
<intersection>327.5 0</intersection>
<intersection>329 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>329,-70,329,-69</points>
<connection>
<GID>391</GID>
<name>IN_B_3</name></connection>
<intersection>-69 3</intersection></vsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323,-82.5,323,-82.5</points>
<connection>
<GID>393</GID>
<name>N_in0</name></connection>
<connection>
<GID>394</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321,-82.5,321,-82.5</points>
<connection>
<GID>394</GID>
<name>N_in0</name></connection>
<connection>
<GID>395</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319,-82.5,319,-82.5</points>
<connection>
<GID>395</GID>
<name>N_in0</name></connection>
<connection>
<GID>396</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325.5,-81.5,325.5,-78</points>
<connection>
<GID>391</GID>
<name>OUT_3</name></connection>
<intersection>-81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>325.5,-81.5,330.5,-81.5</points>
<connection>
<GID>392</GID>
<name>IN_3</name></connection>
<intersection>325.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326.5,-82.5,326.5,-78</points>
<connection>
<GID>391</GID>
<name>OUT_2</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>326.5,-82.5,330.5,-82.5</points>
<connection>
<GID>392</GID>
<name>IN_2</name></connection>
<intersection>326.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327.5,-83.5,327.5,-78</points>
<connection>
<GID>391</GID>
<name>OUT_1</name></connection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>327.5,-83.5,330.5,-83.5</points>
<connection>
<GID>392</GID>
<name>IN_1</name></connection>
<intersection>327.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328.5,-84.5,328.5,-78</points>
<connection>
<GID>391</GID>
<name>OUT_0</name></connection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>328.5,-84.5,330.5,-84.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>328.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-60,337,-57</points>
<connection>
<GID>390</GID>
<name>IN_1</name></connection>
<connection>
<GID>297</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,-60,333,-58</points>
<connection>
<GID>389</GID>
<name>IN_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>336,-58,336,-57</points>
<connection>
<GID>297</GID>
<name>OUT_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>333,-58,336,-58</points>
<intersection>333 0</intersection>
<intersection>336 1</intersection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329,-60,329,-58</points>
<connection>
<GID>388</GID>
<name>IN_1</name></connection>
<intersection>-58 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>335,-58,335,-57</points>
<connection>
<GID>297</GID>
<name>OUT_2</name></connection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>329,-58,335,-58</points>
<intersection>329 0</intersection>
<intersection>335 1</intersection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,-57.5,334,-57</points>
<connection>
<GID>297</GID>
<name>OUT_3</name></connection>
<intersection>-57.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>325,-60,325,-57.5</points>
<connection>
<GID>387</GID>
<name>IN_1</name></connection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>325,-57.5,334,-57.5</points>
<intersection>325 1</intersection>
<intersection>334 0</intersection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326,-40,326,-40</points>
<connection>
<GID>398</GID>
<name>OUT</name></connection>
<connection>
<GID>290</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325,-34,325,-34</points>
<connection>
<GID>398</GID>
<name>IN_1</name></connection>
<connection>
<GID>399</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>574,-38.5,574,25</points>
<intersection>-38.5 1</intersection>
<intersection>25 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>530,-38.5,584,-38.5</points>
<connection>
<GID>310</GID>
<name>IN_2</name></connection>
<intersection>530 6</intersection>
<intersection>574 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>530,-38.5,530,-23</points>
<connection>
<GID>311</GID>
<name>IN_2</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>553.5,25,574,25</points>
<connection>
<GID>411</GID>
<name>OUT_2</name></connection>
<intersection>574 0</intersection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350,-46.5,351.5,-46.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<connection>
<GID>284</GID>
<name>A_less_B</name></connection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>343.5,-52,359,-52</points>
<connection>
<GID>288</GID>
<name>carry_out</name></connection>
<intersection>343.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>343.5,-52,343.5,-38.5</points>
<connection>
<GID>297</GID>
<name>carry_in</name></connection>
<intersection>-52 1</intersection>
<intersection>-38.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>329,-38.5,343.5,-38.5</points>
<intersection>329 5</intersection>
<intersection>343.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>329,-38.5,329,-34</points>
<intersection>-38.5 4</intersection>
<intersection>-34 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>327,-34,329,-34</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>329 5</intersection></hsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>575.5,-39.5,575.5,26</points>
<intersection>-39.5 1</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>528,-39.5,584,-39.5</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<intersection>528 8</intersection>
<intersection>575.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>553.5,26,575.5,26</points>
<connection>
<GID>411</GID>
<name>OUT_1</name></connection>
<intersection>575.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>528,-39.5,528,-24</points>
<intersection>-39.5 1</intersection>
<intersection>-24 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>528,-24,530,-24</points>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<intersection>528 8</intersection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>577,-40.5,577,27</points>
<intersection>-40.5 1</intersection>
<intersection>27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525.5,-40.5,584,-40.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>525.5 7</intersection>
<intersection>577 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>553.5,27,577,27</points>
<connection>
<GID>411</GID>
<name>OUT_0</name></connection>
<intersection>577 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>525.5,-40.5,525.5,-25</points>
<intersection>-40.5 1</intersection>
<intersection>-25 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>525.5,-25,530,-25</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>525.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>548.5,11.5,548.5,17.5</points>
<connection>
<GID>412</GID>
<name>carry_in</name></connection>
<connection>
<GID>411</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515,-32.5,515,5</points>
<connection>
<GID>673</GID>
<name>OUT_0</name></connection>
<intersection>-28.5 16</intersection>
<intersection>-12 6</intersection>
<intersection>5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>510,5,516,5</points>
<connection>
<GID>313</GID>
<name>clear</name></connection>
<intersection>515 0</intersection>
<intersection>516 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>510,-12,515,-12</points>
<intersection>510 13</intersection>
<intersection>515 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>516,5,516,22</points>
<intersection>5 5</intersection>
<intersection>22 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>511,22,516,22</points>
<connection>
<GID>312</GID>
<name>clear</name></connection>
<intersection>516 7</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>510,-12,510,-11</points>
<connection>
<GID>325</GID>
<name>clear</name></connection>
<intersection>-12 6</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>515,-28.5,535,-28.5</points>
<intersection>515 0</intersection>
<intersection>535 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>535,-28.5,535,-27</points>
<connection>
<GID>311</GID>
<name>clear</name></connection>
<intersection>-28.5 16</intersection></vsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>501,24.5,501,28.5</points>
<intersection>24.5 2</intersection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>501,28.5,507.5,28.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>501 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>495,24.5,501,24.5</points>
<connection>
<GID>223</GID>
<name>OUT_3</name></connection>
<intersection>501 0</intersection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502,22.5,502,27.5</points>
<intersection>22.5 2</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>502,27.5,507.5,27.5</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<intersection>502 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>495,22.5,502,22.5</points>
<connection>
<GID>223</GID>
<name>OUT_2</name></connection>
<intersection>502 0</intersection></hsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502,20.5,502,26.5</points>
<intersection>20.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>495,20.5,502,20.5</points>
<connection>
<GID>223</GID>
<name>OUT_1</name></connection>
<intersection>502 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>502,26.5,507.5,26.5</points>
<connection>
<GID>312</GID>
<name>IN_2</name></connection>
<intersection>502 0</intersection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>503.5,18.5,503.5,25.5</points>
<intersection>18.5 1</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>495,18.5,503.5,18.5</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>503.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503.5,25.5,507.5,25.5</points>
<connection>
<GID>312</GID>
<name>IN_3</name></connection>
<intersection>503.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>501,8,501,8.5</points>
<intersection>8 2</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>501,8.5,506.5,8.5</points>
<connection>
<GID>313</GID>
<name>IN_3</name></connection>
<intersection>501 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>494.5,8,501,8</points>
<connection>
<GID>260</GID>
<name>OUT_3</name></connection>
<intersection>501 0</intersection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502,6,502,9.5</points>
<intersection>6 2</intersection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>502,9.5,506.5,9.5</points>
<connection>
<GID>313</GID>
<name>IN_2</name></connection>
<intersection>502 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>494.5,6,502,6</points>
<connection>
<GID>260</GID>
<name>OUT_2</name></connection>
<intersection>502 0</intersection></hsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>503,4,503,10.5</points>
<intersection>4 2</intersection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503,10.5,506.5,10.5</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>503 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>494.5,4,503,4</points>
<connection>
<GID>260</GID>
<name>OUT_1</name></connection>
<intersection>503 0</intersection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>498.5,2,498.5,14</points>
<intersection>2 2</intersection>
<intersection>14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>498.5,14,506.5,14</points>
<intersection>498.5 0</intersection>
<intersection>506.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>494.5,2,498.5,2</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<intersection>498.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>506.5,11.5,506.5,14</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>14 1</intersection></vsegment></shape></wire>
<wire>
<ID>768</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,15,510,15.5</points>
<connection>
<GID>313</GID>
<name>shift_enable</name></connection>
<intersection>15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>509.5,15.5,509.5,16</points>
<connection>
<GID>383</GID>
<name>OUT_0</name></connection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>509.5,15.5,510,15.5</points>
<intersection>509.5 1</intersection>
<intersection>510 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-22.5313,2747.87,1201.47,2142.87</PageViewport></page 3>
<page 4>
<PageViewport>365.559,2045.3,858.485,1801.65</PageViewport>
<gate>
<ID>585</ID>
<type>DD_KEYPAD_HEX</type>
<position>491.5,1937</position>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>414</ID>
<type>DA_FROM</type>
<position>406.5,1963</position>
<input>
<ID>IN_0</ID>603 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i1</lparam></gate>
<gate>
<ID>417</ID>
<type>DA_FROM</type>
<position>406.5,1965</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i2</lparam></gate>
<gate>
<ID>422</ID>
<type>DA_FROM</type>
<position>406.5,1967</position>
<input>
<ID>IN_0</ID>604 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i3</lparam></gate>
<gate>
<ID>424</ID>
<type>DA_FROM</type>
<position>406.5,1969</position>
<input>
<ID>IN_0</ID>622 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i4</lparam></gate>
<gate>
<ID>425</ID>
<type>DA_FROM</type>
<position>406.5,1971</position>
<input>
<ID>IN_0</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i5</lparam></gate>
<gate>
<ID>427</ID>
<type>DA_FROM</type>
<position>406.5,1973</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i6</lparam></gate>
<gate>
<ID>430</ID>
<type>DA_FROM</type>
<position>406.5,1975</position>
<input>
<ID>IN_0</ID>606 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i7</lparam></gate>
<gate>
<ID>431</ID>
<type>DA_FROM</type>
<position>406.5,1977</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i8</lparam></gate>
<gate>
<ID>432</ID>
<type>DA_FROM</type>
<position>406.5,1979</position>
<input>
<ID>IN_0</ID>612 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i9</lparam></gate>
<gate>
<ID>433</ID>
<type>AE_REGISTER8</type>
<position>441,1962.5</position>
<input>
<ID>IN_0</ID>628 </input>
<input>
<ID>IN_1</ID>627 </input>
<input>
<ID>IN_2</ID>626 </input>
<input>
<ID>IN_3</ID>625 </input>
<output>
<ID>OUT_0</ID>716 </output>
<output>
<ID>OUT_1</ID>717 </output>
<output>
<ID>OUT_2</ID>718 </output>
<output>
<ID>OUT_3</ID>719 </output>
<input>
<ID>clock</ID>738 </input>
<input>
<ID>load</ID>738 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>434</ID>
<type>AE_OR2</type>
<position>461,1934</position>
<input>
<ID>IN_0</ID>746 </input>
<input>
<ID>IN_1</ID>745 </input>
<output>
<ID>OUT</ID>744 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>435</ID>
<type>DA_FROM</type>
<position>460,1929</position>
<input>
<ID>IN_0</ID>746 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID +</lparam></gate>
<gate>
<ID>436</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>433,1970</position>
<input>
<ID>IN_0</ID>615 </input>
<input>
<ID>IN_1</ID>616 </input>
<input>
<ID>IN_2</ID>620 </input>
<input>
<ID>IN_3</ID>619 </input>
<output>
<ID>OUT_0</ID>628 </output>
<output>
<ID>OUT_1</ID>627 </output>
<output>
<ID>OUT_2</ID>626 </output>
<output>
<ID>OUT_3</ID>625 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>437</ID>
<type>DE_OR8</type>
<position>422,1959</position>
<input>
<ID>IN_0</ID>614 </input>
<input>
<ID>IN_1</ID>614 </input>
<input>
<ID>IN_2</ID>614 </input>
<input>
<ID>IN_3</ID>612 </input>
<input>
<ID>IN_4</ID>603 </input>
<input>
<ID>IN_5</ID>604 </input>
<input>
<ID>IN_6</ID>605 </input>
<input>
<ID>IN_7</ID>606 </input>
<output>
<ID>OUT</ID>615 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>438</ID>
<type>FF_GND</type>
<position>418,1960.5</position>
<output>
<ID>OUT_0</ID>614 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>439</ID>
<type>AE_OR2</type>
<position>422,1981</position>
<input>
<ID>IN_0</ID>612 </input>
<input>
<ID>IN_1</ID>621 </input>
<output>
<ID>OUT</ID>619 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>440</ID>
<type>AE_OR4</type>
<position>421,1967</position>
<input>
<ID>IN_0</ID>606 </input>
<input>
<ID>IN_1</ID>618 </input>
<input>
<ID>IN_2</ID>604 </input>
<input>
<ID>IN_3</ID>617 </input>
<output>
<ID>OUT</ID>616 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>441</ID>
<type>AE_OR4</type>
<position>421,1975</position>
<input>
<ID>IN_0</ID>606 </input>
<input>
<ID>IN_1</ID>618 </input>
<input>
<ID>IN_2</ID>605 </input>
<input>
<ID>IN_3</ID>622 </input>
<output>
<ID>OUT</ID>620 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>444</ID>
<type>DA_FROM</type>
<position>406.5,1961</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID i0</lparam></gate>
<gate>
<ID>471</ID>
<type>AE_OR4</type>
<position>430,1959</position>
<input>
<ID>IN_0</ID>619 </input>
<input>
<ID>IN_1</ID>620 </input>
<input>
<ID>IN_2</ID>616 </input>
<input>
<ID>IN_3</ID>615 </input>
<output>
<ID>OUT</ID>623 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>472</ID>
<type>AE_OR2</type>
<position>437,1955.5</position>
<input>
<ID>IN_0</ID>623 </input>
<input>
<ID>IN_1</ID>624 </input>
<output>
<ID>OUT</ID>738 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>475</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>461,1962</position>
<input>
<ID>IN_0</ID>716 </input>
<input>
<ID>IN_1</ID>717 </input>
<input>
<ID>IN_2</ID>718 </input>
<input>
<ID>IN_3</ID>719 </input>
<output>
<ID>carry_out</ID>700 </output>
<input>
<ID>clear</ID>744 </input>
<input>
<ID>clock</ID>741 </input>
<input>
<ID>load</ID>598 </input>
<input>
<ID>shift_enable</ID>701 </input>
<input>
<ID>shift_left</ID>720 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>476</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>461,1949</position>
<input>
<ID>carry_in</ID>700 </input>
<input>
<ID>clear</ID>744 </input>
<input>
<ID>clock</ID>741 </input>
<input>
<ID>shift_enable</ID>701 </input>
<input>
<ID>shift_left</ID>739 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>477</ID>
<type>BB_CLOCK</type>
<position>406,1939</position>
<output>
<ID>CLK</ID>709 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>478</ID>
<type>BA_SHIFT_REGISTER_4</type>
<position>414,1945.5</position>
<input>
<ID>IN_0</ID>710 </input>
<output>
<ID>OUT_0</ID>711 </output>
<output>
<ID>OUT_1</ID>712 </output>
<output>
<ID>OUT_2</ID>713 </output>
<output>
<ID>OUT_3</ID>714 </output>
<output>
<ID>carry_out</ID>737 </output>
<input>
<ID>clear</ID>737 </input>
<input>
<ID>clock</ID>709 </input>
<input>
<ID>load</ID>738 </input>
<input>
<ID>shift_enable</ID>710 </input>
<input>
<ID>shift_left</ID>710 </input>
<gparam>VALUE_BOX -0.8,-1.3,0.8,1.3</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>479</ID>
<type>EE_VDD</type>
<position>409.5,1947</position>
<output>
<ID>OUT_0</ID>710 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>480</ID>
<type>AE_OR4</type>
<position>422.5,1945.5</position>
<input>
<ID>IN_0</ID>711 </input>
<input>
<ID>IN_1</ID>712 </input>
<input>
<ID>IN_2</ID>713 </input>
<input>
<ID>IN_3</ID>714 </input>
<output>
<ID>OUT</ID>721 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>289</ID>
<type>AE_SMALL_INVERTER</type>
<position>451.5,1941.5</position>
<input>
<ID>IN_0</ID>599 </input>
<output>
<ID>OUT_0</ID>598 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>485</ID>
<type>GA_LED</type>
<position>435.5,1944.5</position>
<input>
<ID>N_in0</ID>735 </input>
<input>
<ID>N_in1</ID>715 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>AE_SMALL_INVERTER</type>
<position>439.5,1941.5</position>
<input>
<ID>IN_0</ID>601 </input>
<output>
<ID>OUT_0</ID>600 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>491</ID>
<type>DE_TO</type>
<position>438.5,1944.5</position>
<input>
<ID>IN_0</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cc</lparam></gate>
<gate>
<ID>492</ID>
<type>EE_VDD</type>
<position>463,1968</position>
<output>
<ID>OUT_0</ID>720 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>493</ID>
<type>EE_VDD</type>
<position>464,1956</position>
<output>
<ID>OUT_0</ID>739 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>494</ID>
<type>AA_AND2</type>
<position>431.5,1944.5</position>
<input>
<ID>IN_0</ID>721 </input>
<input>
<ID>IN_1</ID>736 </input>
<output>
<ID>OUT</ID>735 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>495</ID>
<type>AE_SMALL_INVERTER</type>
<position>418,1939</position>
<input>
<ID>IN_0</ID>709 </input>
<output>
<ID>OUT_0</ID>596 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>303</ID>
<type>AE_SMALL_INVERTER</type>
<position>443.5,1941.5</position>
<input>
<ID>IN_0</ID>600 </input>
<output>
<ID>OUT_0</ID>602 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>496</ID>
<type>AE_SMALL_INVERTER</type>
<position>422,1939</position>
<input>
<ID>IN_0</ID>596 </input>
<output>
<ID>OUT_0</ID>736 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>497</ID>
<type>DA_FROM</type>
<position>461,1973</position>
<input>
<ID>IN_0</ID>701 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID cc</lparam></gate>
<gate>
<ID>498</ID>
<type>AE_SMALL_INVERTER</type>
<position>439.5,1939</position>
<input>
<ID>IN_0</ID>736 </input>
<output>
<ID>OUT_0</ID>740 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>499</ID>
<type>AE_SMALL_INVERTER</type>
<position>443.5,1939</position>
<input>
<ID>IN_0</ID>740 </input>
<output>
<ID>OUT_0</ID>743 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>500</ID>
<type>AE_SMALL_INVERTER</type>
<position>447.5,1939</position>
<input>
<ID>IN_0</ID>743 </input>
<output>
<ID>OUT_0</ID>742 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>501</ID>
<type>AE_SMALL_INVERTER</type>
<position>451.5,1939</position>
<input>
<ID>IN_0</ID>742 </input>
<output>
<ID>OUT_0</ID>741 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>503</ID>
<type>CC_PULSE</type>
<position>399.5,1979.5</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>505</ID>
<type>CC_PULSE</type>
<position>399.5,1976.5</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>507</ID>
<type>CC_PULSE</type>
<position>399.5,1974</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>509</ID>
<type>CC_PULSE</type>
<position>399.5,1971.5</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>511</ID>
<type>CC_PULSE</type>
<position>399.5,1969</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>513</ID>
<type>CC_PULSE</type>
<position>399.5,1966.5</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>515</ID>
<type>CC_PULSE</type>
<position>399.5,1964</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>517</ID>
<type>CC_PULSE</type>
<position>399.5,1961</position>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>327</ID>
<type>DA_FROM</type>
<position>462,1929</position>
<input>
<ID>IN_0</ID>745 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>328</ID>
<type>DE_TO</type>
<position>447.5,1950</position>
<input>
<ID>IN_0</ID>738 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID klaw</lparam></gate>
<gate>
<ID>521</ID>
<type>DD_KEYPAD_HEX</type>
<position>491.5,1949.5</position>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>522</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>510.5,1967.5</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>166</ID>
<type>AE_SMALL_INVERTER</type>
<position>431.5,1941.5</position>
<input>
<ID>IN_0</ID>714 </input>
<output>
<ID>OUT_0</ID>597 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>167</ID>
<type>AE_SMALL_INVERTER</type>
<position>435.5,1941.5</position>
<input>
<ID>IN_0</ID>597 </input>
<output>
<ID>OUT_0</ID>601 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>168</ID>
<type>AE_SMALL_INVERTER</type>
<position>447.5,1941.5</position>
<input>
<ID>IN_0</ID>602 </input>
<output>
<ID>OUT_0</ID>599 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>560</ID>
<type>AE_REGISTER8</type>
<position>497.5,1962.5</position>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>420,1939,420,1939</points>
<connection>
<GID>495</GID>
<name>OUT_0</name></connection>
<connection>
<GID>496</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>433.5,1941.5,433.5,1941.5</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<connection>
<GID>167</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,1941.5,455.5,1969.5</points>
<intersection>1941.5 1</intersection>
<intersection>1969.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>453.5,1941.5,455.5,1941.5</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<intersection>455.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>455.5,1969.5,462,1969.5</points>
<intersection>455.5 0</intersection>
<intersection>462 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>462,1967,462,1969.5</points>
<connection>
<GID>475</GID>
<name>load</name></connection>
<intersection>1969.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449.5,1941.5,449.5,1941.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>441.5,1941.5,441.5,1941.5</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<connection>
<GID>303</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437.5,1941.5,437.5,1941.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445.5,1941.5,445.5,1941.5</points>
<connection>
<GID>303</GID>
<name>OUT_0</name></connection>
<connection>
<GID>168</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>412.5,1955.5,412.5,1963</points>
<intersection>1955.5 2</intersection>
<intersection>1963 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1963,412.5,1963</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>412.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>412.5,1955.5,419,1955.5</points>
<connection>
<GID>437</GID>
<name>IN_4</name></connection>
<intersection>412.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413,1956.5,413,1967</points>
<intersection>1956.5 2</intersection>
<intersection>1966 3</intersection>
<intersection>1967 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1967,413,1967</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413,1956.5,419,1956.5</points>
<connection>
<GID>437</GID>
<name>IN_5</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>413,1966,418,1966</points>
<connection>
<GID>440</GID>
<name>IN_2</name></connection>
<intersection>413 0</intersection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413.5,1957.5,413.5,1974</points>
<intersection>1957.5 2</intersection>
<intersection>1971 1</intersection>
<intersection>1974 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1971,413.5,1971</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>413.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413.5,1957.5,419,1957.5</points>
<connection>
<GID>437</GID>
<name>IN_6</name></connection>
<intersection>413.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>413.5,1974,418,1974</points>
<connection>
<GID>441</GID>
<name>IN_2</name></connection>
<intersection>413.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>414,1958.5,414,1978</points>
<intersection>1958.5 2</intersection>
<intersection>1970 3</intersection>
<intersection>1975 1</intersection>
<intersection>1978 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1975,414,1975</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>414 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>414,1958.5,419,1958.5</points>
<connection>
<GID>437</GID>
<name>IN_7</name></connection>
<intersection>414 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>414,1970,418,1970</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>414 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>414,1978,418,1978</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>414 0</intersection></hsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>414.5,1959.5,414.5,1982</points>
<intersection>1959.5 2</intersection>
<intersection>1979 1</intersection>
<intersection>1982 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1979,414.5,1979</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<intersection>414.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>414.5,1959.5,419,1959.5</points>
<connection>
<GID>437</GID>
<name>IN_3</name></connection>
<intersection>414.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>414.5,1982,419,1982</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<intersection>414.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>419,1960.5,419,1962.5</points>
<connection>
<GID>438</GID>
<name>OUT_0</name></connection>
<connection>
<GID>437</GID>
<name>IN_2</name></connection>
<connection>
<GID>437</GID>
<name>IN_1</name></connection>
<connection>
<GID>437</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426,1956,426,1969</points>
<connection>
<GID>437</GID>
<name>OUT</name></connection>
<intersection>1956 6</intersection>
<intersection>1969 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>426,1969,430,1969</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<intersection>426 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>426,1956,427,1956</points>
<connection>
<GID>471</GID>
<name>IN_3</name></connection>
<intersection>426 0</intersection></hsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,1958,425.5,1970</points>
<intersection>1958 3</intersection>
<intersection>1967 2</intersection>
<intersection>1970 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425.5,1970,430,1970</points>
<connection>
<GID>436</GID>
<name>IN_1</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>425,1967,425.5,1967</points>
<connection>
<GID>440</GID>
<name>OUT</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>425.5,1958,427,1958</points>
<connection>
<GID>471</GID>
<name>IN_2</name></connection>
<intersection>425.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413,1964,413,1965</points>
<intersection>1964 2</intersection>
<intersection>1965 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1965,413,1965</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413,1964,418,1964</points>
<connection>
<GID>440</GID>
<name>IN_3</name></connection>
<intersection>413 0</intersection></hsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413,1968,413,1976</points>
<intersection>1968 2</intersection>
<intersection>1973 1</intersection>
<intersection>1976 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1973,413,1973</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413,1968,418,1968</points>
<connection>
<GID>440</GID>
<name>IN_1</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>413,1976,418,1976</points>
<connection>
<GID>441</GID>
<name>IN_1</name></connection>
<intersection>413 0</intersection></hsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426,1972,426,1981</points>
<intersection>1972 3</intersection>
<intersection>1981 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>425,1981,426,1981</points>
<connection>
<GID>439</GID>
<name>OUT</name></connection>
<intersection>426 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>426,1972,430,1972</points>
<connection>
<GID>436</GID>
<name>IN_3</name></connection>
<intersection>426 0</intersection>
<intersection>427 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>427,1962,427,1972</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<intersection>1972 3</intersection></vsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,1971,425.5,1975</points>
<intersection>1971 1</intersection>
<intersection>1975 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425.5,1971,430,1971</points>
<connection>
<GID>436</GID>
<name>IN_2</name></connection>
<intersection>425.5 0</intersection>
<intersection>426.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>425,1975,425.5,1975</points>
<connection>
<GID>441</GID>
<name>OUT</name></connection>
<intersection>425.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>426.5,1960,426.5,1971</points>
<intersection>1960 6</intersection>
<intersection>1971 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>426.5,1960,427,1960</points>
<connection>
<GID>471</GID>
<name>IN_1</name></connection>
<intersection>426.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413.5,1977,413.5,1980</points>
<intersection>1977 1</intersection>
<intersection>1980 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1977,413.5,1977</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<intersection>413.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413.5,1980,419,1980</points>
<connection>
<GID>439</GID>
<name>IN_1</name></connection>
<intersection>413.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413,1969,413,1972</points>
<intersection>1969 1</intersection>
<intersection>1972 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1969,413,1969</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>413 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413,1972,418,1972</points>
<connection>
<GID>441</GID>
<name>IN_3</name></connection>
<intersection>413 0</intersection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>434,1956.5,434,1959</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<connection>
<GID>471</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>412,1954.5,412,1961</points>
<intersection>1954.5 2</intersection>
<intersection>1961 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,1961,412,1961</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>412 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>412,1954.5,434,1954.5</points>
<connection>
<GID>472</GID>
<name>IN_1</name></connection>
<intersection>412 0</intersection></hsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431.5,1962.5,431.5,1966</points>
<connection>
<GID>436</GID>
<name>OUT_3</name></connection>
<intersection>1962.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>431.5,1962.5,437,1962.5</points>
<connection>
<GID>433</GID>
<name>IN_3</name></connection>
<intersection>431.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432.5,1961.5,432.5,1966</points>
<connection>
<GID>436</GID>
<name>OUT_2</name></connection>
<intersection>1961.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,1961.5,437,1961.5</points>
<connection>
<GID>433</GID>
<name>IN_2</name></connection>
<intersection>432.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>433.5,1960.5,433.5,1966</points>
<connection>
<GID>436</GID>
<name>OUT_1</name></connection>
<intersection>1960.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>433.5,1960.5,437,1960.5</points>
<connection>
<GID>433</GID>
<name>IN_1</name></connection>
<intersection>433.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,1959.5,434.5,1966</points>
<connection>
<GID>436</GID>
<name>OUT_0</name></connection>
<intersection>1959.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,1959.5,437,1959.5</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<vsegment>
<ID>20</ID>
<points>459.5,1954,459.5,1957</points>
<connection>
<GID>476</GID>
<name>carry_in</name></connection>
<connection>
<GID>475</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>466,1954.5,466,1971</points>
<intersection>1954.5 20</intersection>
<intersection>1971 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>461,1971,466,1971</points>
<intersection>461 22</intersection>
<intersection>466 1</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>461,1954.5,466,1954.5</points>
<intersection>461 21</intersection>
<intersection>466 1</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>461,1954,461,1954.5</points>
<connection>
<GID>476</GID>
<name>shift_enable</name></connection>
<intersection>1954.5 20</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>461,1967,461,1971</points>
<connection>
<GID>475</GID>
<name>shift_enable</name></connection>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<intersection>1971 18</intersection></vsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<vsegment>
<ID>18</ID>
<points>415,1939,415,1940.5</points>
<connection>
<GID>478</GID>
<name>clock</name></connection>
<intersection>1939 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>410,1939,416,1939</points>
<connection>
<GID>477</GID>
<name>CLK</name></connection>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>415 18</intersection></hsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>410.5,1947,410.5,1951.5</points>
<connection>
<GID>479</GID>
<name>OUT_0</name></connection>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>1951.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>410.5,1951.5,416,1951.5</points>
<intersection>410.5 0</intersection>
<intersection>414 14</intersection>
<intersection>416 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>416,1950.5,416,1951.5</points>
<connection>
<GID>478</GID>
<name>shift_left</name></connection>
<intersection>1951.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>414,1950.5,414,1951.5</points>
<connection>
<GID>478</GID>
<name>shift_enable</name></connection>
<intersection>1951.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>418,1947,418,1948.5</points>
<intersection>1947 1</intersection>
<intersection>1948.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>417.5,1947,418,1947</points>
<connection>
<GID>478</GID>
<name>OUT_0</name></connection>
<intersection>418 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>418,1948.5,419.5,1948.5</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>418 0</intersection></hsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>417.5,1946.5,419.5,1946.5</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>417.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>417.5,1946,417.5,1946.5</points>
<connection>
<GID>478</GID>
<name>OUT_1</name></connection>
<intersection>1946.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>417.5,1944.5,419.5,1944.5</points>
<connection>
<GID>480</GID>
<name>IN_2</name></connection>
<intersection>417.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>417.5,1944.5,417.5,1945</points>
<connection>
<GID>478</GID>
<name>OUT_2</name></connection>
<intersection>1944.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>417.5,1941.5,417.5,1944</points>
<connection>
<GID>478</GID>
<name>OUT_3</name></connection>
<intersection>1941.5 12</intersection>
<intersection>1942.5 15</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>417.5,1941.5,429.5,1941.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>417.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>417.5,1942.5,419.5,1942.5</points>
<connection>
<GID>480</GID>
<name>IN_3</name></connection>
<intersection>417.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436.5,1944.5,436.5,1944.5</points>
<connection>
<GID>485</GID>
<name>N_in1</name></connection>
<connection>
<GID>491</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>453,1959.5,453,1963.5</points>
<intersection>1959.5 1</intersection>
<intersection>1963.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445,1959.5,453,1959.5</points>
<connection>
<GID>433</GID>
<name>OUT_0</name></connection>
<intersection>453 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>453,1963.5,457.5,1963.5</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>453 0</intersection></hsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448.5,1960.5,448.5,1963</points>
<intersection>1960.5 1</intersection>
<intersection>1963 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445,1960.5,448.5,1960.5</points>
<connection>
<GID>433</GID>
<name>OUT_1</name></connection>
<intersection>448.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448.5,1963,457.5,1963</points>
<intersection>448.5 0</intersection>
<intersection>457.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>457.5,1962.5,457.5,1963</points>
<connection>
<GID>475</GID>
<name>IN_1</name></connection>
<intersection>1963 2</intersection></vsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>445,1961.5,457.5,1961.5</points>
<connection>
<GID>433</GID>
<name>OUT_2</name></connection>
<connection>
<GID>475</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450,1960.5,450,1962.5</points>
<intersection>1960.5 2</intersection>
<intersection>1962.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445,1962.5,450,1962.5</points>
<connection>
<GID>433</GID>
<name>OUT_3</name></connection>
<intersection>450 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450,1960.5,457.5,1960.5</points>
<connection>
<GID>475</GID>
<name>IN_3</name></connection>
<intersection>450 0</intersection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>463,1967,463,1967</points>
<connection>
<GID>475</GID>
<name>shift_left</name></connection>
<connection>
<GID>492</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>426.5,1945.5,428.5,1945.5</points>
<connection>
<GID>480</GID>
<name>OUT</name></connection>
<connection>
<GID>494</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,1944.5,434.5,1944.5</points>
<connection>
<GID>485</GID>
<name>N_in0</name></connection>
<connection>
<GID>494</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428,1939,428,1943.5</points>
<intersection>1939 5</intersection>
<intersection>1943.5 15</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>424,1939,437.5,1939</points>
<connection>
<GID>496</GID>
<name>OUT_0</name></connection>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>428 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>428,1943.5,428.5,1943.5</points>
<connection>
<GID>494</GID>
<name>IN_1</name></connection>
<intersection>428 0</intersection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412.5,1940.5,414,1940.5</points>
<connection>
<GID>478</GID>
<name>clear</name></connection>
<connection>
<GID>478</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>415,1950.5,415,1953</points>
<connection>
<GID>478</GID>
<name>load</name></connection>
<intersection>1953 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>415,1953,447,1953</points>
<intersection>415 0</intersection>
<intersection>445.5 16</intersection>
<intersection>447 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>447,1953,447,1973</points>
<intersection>1953 1</intersection>
<intersection>1955.5 5</intersection>
<intersection>1973 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>440,1973,447,1973</points>
<intersection>440 7</intersection>
<intersection>447 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>440,1955.5,447,1955.5</points>
<connection>
<GID>472</GID>
<name>OUT</name></connection>
<intersection>440 8</intersection>
<intersection>447 2</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>440,1968.5,440,1973</points>
<connection>
<GID>433</GID>
<name>load</name></connection>
<intersection>1973 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>440,1955.5,440,1957.5</points>
<connection>
<GID>433</GID>
<name>clock</name></connection>
<intersection>1955.5 5</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>445.5,1950,445.5,1953</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>1953 1</intersection></vsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>463,1954,463,1956</points>
<connection>
<GID>493</GID>
<name>OUT_0</name></connection>
<connection>
<GID>476</GID>
<name>shift_left</name></connection></vsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>441.5,1939,441.5,1939</points>
<connection>
<GID>498</GID>
<name>OUT_0</name></connection>
<connection>
<GID>499</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>465,1939,465,1957</points>
<intersection>1939 8</intersection>
<intersection>1944 5</intersection>
<intersection>1957 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>462,1944,465,1944</points>
<connection>
<GID>476</GID>
<name>clock</name></connection>
<intersection>465 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>462,1957,465,1957</points>
<connection>
<GID>475</GID>
<name>clock</name></connection>
<intersection>465 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>453.5,1939,465,1939</points>
<connection>
<GID>501</GID>
<name>OUT_0</name></connection>
<intersection>465 0</intersection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449.5,1939,449.5,1939</points>
<connection>
<GID>500</GID>
<name>OUT_0</name></connection>
<connection>
<GID>501</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445.5,1939,445.5,1939</points>
<connection>
<GID>499</GID>
<name>OUT_0</name></connection>
<connection>
<GID>500</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>744</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454.5,1940,454.5,1957</points>
<intersection>1940 4</intersection>
<intersection>1957 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>454.5,1957,461,1957</points>
<connection>
<GID>475</GID>
<name>clear</name></connection>
<intersection>454.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>454.5,1940,461,1940</points>
<intersection>454.5 0</intersection>
<intersection>461 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>461,1937,461,1944</points>
<connection>
<GID>434</GID>
<name>OUT</name></connection>
<connection>
<GID>476</GID>
<name>clear</name></connection>
<intersection>1940 4</intersection></vsegment></shape></wire>
<wire>
<ID>745</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>462,1931,462,1931</points>
<connection>
<GID>434</GID>
<name>IN_1</name></connection>
<connection>
<GID>327</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>746</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>460,1931,460,1931</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<connection>
<GID>435</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-22.5313,2747.87,1201.47,2142.87</PageViewport></page 5>
<page 6>
<PageViewport>-22.5313,2747.87,1201.47,2142.87</PageViewport></page 6>
<page 7>
<PageViewport>-22.5313,2747.87,1201.47,2142.87</PageViewport></page 7>
<page 8>
<PageViewport>-22.5313,2747.87,1201.47,2142.87</PageViewport></page 8>
<page 9>
<PageViewport>-22.5313,2747.87,1201.47,2142.87</PageViewport></page 9></circuit>