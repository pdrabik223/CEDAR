<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-61.5086,-49.2939,153.163,-290.799</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>39,-168.5</position>
<gparam>LABEL_TEXT Zadanie 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>35.5,-10.5</position>
<gparam>LABEL_TEXT Uklad sumy i roznicy zupelnej</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>22.5,-175</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>18.5,-16</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>22.5,-180.5</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>18.5,-21</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>22.5,-185</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>18.5,-26</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>18,-175</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AE_SMALL_INVERTER</type>
<position>28.5,-16</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_SMALL_INVERTER</type>
<position>28.5,-21</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>28.5,-26</position>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>18,-180</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>BA_NAND3</type>
<position>40.5,-17</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>18 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>15</ID>
<type>BA_NAND3</type>
<position>40.5,-23.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>4 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>BA_NAND3</type>
<position>40.5,-30</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>4 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>17.5,-184.5</position>
<gparam>LABEL_TEXT Bi</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>BA_NAND4</type>
<position>52,-27</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>9 </input>
<input>
<ID>IN_3</ID>49 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND2</type>
<position>41,-176</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>57,-27</position>
<input>
<ID>N_in0</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>35,-45</position>
<gparam>LABEL_TEXT Uklad sumy i roznicy zbudowany z XOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>17.5,-50</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>17.5,-56</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>17.5,-61</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_SMALL_INVERTER</type>
<position>33,-175</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AI_XOR2</type>
<position>30.5,-53</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AI_XOR2</type>
<position>37,-60</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>41,-60</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>15.5,-15.5</position>
<gparam>LABEL_TEXT J</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>15.5,-20.5</position>
<gparam>LABEL_TEXT K</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>16,-25.5</position>
<gparam>LABEL_TEXT L</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>60,-26.5</position>
<gparam>LABEL_TEXT M</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>44,-59.5</position>
<gparam>LABEL_TEXT M</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>15,-60.5</position>
<gparam>LABEL_TEXT L</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>14.5,-55.5</position>
<gparam>LABEL_TEXT K</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>15,-49.5</position>
<gparam>LABEL_TEXT J</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>30,-69</position>
<gparam>LABEL_TEXT C0 dla sumatora pe�nego</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>18.5,-78</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>18.5,-81.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>18.5,-89.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>16,-89</position>
<gparam>LABEL_TEXT Ci</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>16,-81</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>16,-77.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND2</type>
<position>41,-182.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>BA_NAND2</type>
<position>32.5,-79</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>BA_NAND2</type>
<position>32.5,-83.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>BA_NAND2</type>
<position>32.5,-88.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND2</type>
<position>41.5,-188</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>BA_NAND3</type>
<position>45,-83.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>22 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>49,-83.5</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>52.5,-83.5</position>
<gparam>LABEL_TEXT Cio</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>20,-101</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>20,-109</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>20,-122</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>17.5,-121.5</position>
<gparam>LABEL_TEXT Ci</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>17.5,-108.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>17.5,-100.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>BA_NAND2</type>
<position>31.5,-102</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_SMALL_INVERTER</type>
<position>40,-102</position>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>BE_NOR2</type>
<position>48,-106</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>AE_SMALL_INVERTER</type>
<position>57.5,-106</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>69</ID>
<type>AI_XOR2</type>
<position>29,-108.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>BA_NAND2</type>
<position>36.5,-114</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_SMALL_INVERTER</type>
<position>41.5,-114</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>72</ID>
<type>AI_XOR2</type>
<position>35,-121</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>GA_LED</type>
<position>60.5,-106</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>64,-106</position>
<gparam>LABEL_TEXT Cio</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>56.5,-121</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>60,-121</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>33,-95</position>
<gparam>LABEL_TEXT Sumator pelny zbudowany z dwoch polsumatorow X+Y+C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>34,-127.5</position>
<gparam>LABEL_TEXT Dwu bitowy sumator rownolegly</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>60,-182.5</position>
<input>
<ID>N_in0</ID>55 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>14,-137.5</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_TOGGLE</type>
<position>14,-144</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>14,-149.5</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_TOGGLE</type>
<position>14,-155</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>85</ID>
<type>BA_NAND2</type>
<position>31,-138.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>AI_XOR3</type>
<position>56,-182.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>56 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>87</ID>
<type>AI_XOR2</type>
<position>31.5,-144</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>88</ID>
<type>BA_NAND2</type>
<position>31,-150</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>AI_XOR2</type>
<position>31.5,-155.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_SMALL_INVERTER</type>
<position>36,-138.5</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>92</ID>
<type>BA_NAND2</type>
<position>41,-156.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AI_XOR2</type>
<position>42,-162</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>BA_NAND2</type>
<position>52.5,-147</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>GA_LED</type>
<position>61,-144</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>GA_LED</type>
<position>61,-147</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>GA_LED</type>
<position>61,-162</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>11,-137</position>
<gparam>LABEL_TEXT X0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>11,-143.5</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>11,-149</position>
<gparam>LABEL_TEXT X1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>10.5,-154.5</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>66,-161.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>66,-146.5</position>
<gparam>LABEL_TEXT Co1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>66,-143.5</position>
<gparam>LABEL_TEXT So</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>BA_NAND3</type>
<position>40.5,-36.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>18 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-27,56,-27</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<connection>
<GID>21</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-21.5,35,-15</points>
<intersection>-21.5 4</intersection>
<intersection>-16 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-16,35,-16</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-15,37.5,-15</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>35,-21.5,37.5,-21.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-30,34,-17</points>
<intersection>-30 3</intersection>
<intersection>-21 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-17,37.5,-17</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-21,34,-21</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-30,37.5,-30</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-32,33,-25.5</points>
<intersection>-32 1</intersection>
<intersection>-26 2</intersection>
<intersection>-25.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-32,37.5,-32</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-26,33,-26</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-25.5,37.5,-25.5</points>
<connection>
<GID>15</GID>
<name>IN_2</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-16,26.5,-16</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>23 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23,-34.5,23,-16</points>
<intersection>-34.5 12</intersection>
<intersection>-28 4</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>23,-28,37.5,-28</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>23 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>23,-34.5,37.5,-34.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>23 3</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-21,26.5,-21</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-36.5,25,-21</points>
<intersection>-36.5 11</intersection>
<intersection>-23.5 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>25,-23.5,37.5,-23.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>25 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>25,-36.5,37.5,-36.5</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>25 3</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-175,38,-175</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>35 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>35,-187,35,-175</points>
<intersection>-187 8</intersection>
<intersection>-175 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>35,-187,38.5,-187</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>35 7</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-185,33.5,-177</points>
<intersection>-185 1</intersection>
<intersection>-183.5 3</intersection>
<intersection>-177 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-185,33.5,-185</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-177,38,-177</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-183.5,38,-183.5</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-30,46,-28</points>
<intersection>-30 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-28,49,-28</points>
<connection>
<GID>19</GID>
<name>IN_2</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-30,46,-30</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-26,46,-23.5</points>
<intersection>-26 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-26,49,-26</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-23.5,46,-23.5</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-24,48,-17</points>
<intersection>-24 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-24,49,-24</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-17,48,-17</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-61,34,-61</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-56,27.5,-56</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>27.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27.5,-56,27.5,-54</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-56 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-52,27.5,-50</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-50,27.5,-50</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-59,33.5,-53</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-59,34,-59</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-60,40,-60</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<connection>
<GID>30</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-175,31,-175</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-38.5,22,-19</points>
<intersection>-38.5 7</intersection>
<intersection>-26 1</intersection>
<intersection>-19 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-26,26.5,-26</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>22,-19,37.5,-19</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>22,-38.5,37.5,-38.5</points>
<connection>
<GID>105</GID>
<name>IN_2</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-83.5,48,-83.5</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<connection>
<GID>54</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-81.5,38.5,-79</points>
<intersection>-81.5 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-79,38.5,-79</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-81.5,42,-81.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-83.5,42,-83.5</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<connection>
<GID>53</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-88.5,38.5,-85.5</points>
<intersection>-88.5 1</intersection>
<intersection>-85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-88.5,38.5,-88.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-85.5,42,-85.5</points>
<connection>
<GID>53</GID>
<name>IN_2</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-78,29.5,-78</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>23.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>23.5,-87.5,23.5,-78</points>
<intersection>-87.5 5</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>23.5,-87.5,29.5,-87.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>23.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-82.5,25,-80</points>
<intersection>-82.5 2</intersection>
<intersection>-81.5 1</intersection>
<intersection>-80 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-81.5,25,-81.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-82.5,29.5,-82.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>25,-80,29.5,-80</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-89.5,29.5,-89.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>26.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26.5,-89.5,26.5,-84.5</points>
<intersection>-89.5 1</intersection>
<intersection>-84.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>26.5,-84.5,29.5,-84.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>26.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-105,43.5,-102</points>
<intersection>-105 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-102,43.5,-102</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-105,45,-105</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-114,43.5,-107</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-107,45,-107</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51,-106,55.5,-106</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-106,59.5,-106</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<connection>
<GID>73</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-121,55.5,-121</points>
<connection>
<GID>75</GID>
<name>N_in0</name></connection>
<connection>
<GID>72</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-122,32,-122</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>25.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>25.5,-122,25.5,-115</points>
<intersection>-122 1</intersection>
<intersection>-115 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>25.5,-115,33.5,-115</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>25.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-120,32,-108.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>-113 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>32,-113,33.5,-113</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>39.5,-114,39.5,-114</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<connection>
<GID>71</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-102,38,-102</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<connection>
<GID>62</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-107.5,24,-101</points>
<intersection>-107.5 2</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-101,28.5,-101</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-107.5,26,-107.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-109.5,25,-103</points>
<intersection>-109.5 3</intersection>
<intersection>-109 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-109,25,-109</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-103,28.5,-103</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25,-109.5,26,-109.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-156.5,46,-148</points>
<intersection>-156.5 3</intersection>
<intersection>-148 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>44,-156.5,46,-156.5</points>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>46,-148,49.5,-148</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-150,41.5,-146</points>
<intersection>-150 3</intersection>
<intersection>-146 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>34,-150,41.5,-150</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>41.5,-146,49.5,-146</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>34,-138.5,34,-138.5</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<connection>
<GID>91</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-161,37,-155.5</points>
<intersection>-161 5</intersection>
<intersection>-155.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>37,-161,39,-161</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>34.5,-155.5,38,-155.5</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-163,38,-138.5</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<intersection>-163 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>38,-163,39,-163</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>45,-162,60,-162</points>
<connection>
<GID>97</GID>
<name>N_in0</name></connection>
<connection>
<GID>93</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>55.5,-147,60,-147</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<connection>
<GID>96</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>34.5,-144,60,-144</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<connection>
<GID>95</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>16,-137.5,28.5,-137.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>28.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>28.5,-143,28.5,-137.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-137.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-144,21.5,-139.5</points>
<intersection>-144 4</intersection>
<intersection>-139.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>21.5,-139.5,28.5,-139.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection>
<intersection>28.5 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>16,-144,21.5,-144</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>21.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>28.5,-145,28.5,-139.5</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>-139.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-154.5,22,-149.5</points>
<intersection>-154.5 5</intersection>
<intersection>-149.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>22,-154.5,28.5,-154.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection>
<intersection>28 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>16,-149.5,22,-149.5</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>22 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>28,-154.5,28,-149</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>-154.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-156.5,22,-155</points>
<intersection>-156.5 5</intersection>
<intersection>-155 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>22,-156.5,28.5,-156.5</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection>
<intersection>28 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>16,-155,22,-155</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>22 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>28,-156.5,28,-151</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>-156.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-36.5,46,-30</points>
<intersection>-36.5 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-30,49,-30</points>
<connection>
<GID>19</GID>
<name>IN_3</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-36.5,46,-36.5</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-189,31,-180.5</points>
<intersection>-189 4</intersection>
<intersection>-181.5 2</intersection>
<intersection>-180.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-180.5,31,-180.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-181.5,38,-181.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>31,-189,38.5,-189</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-182.5,59,-182.5</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<connection>
<GID>79</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-188,48.5,-184.5</points>
<intersection>-188 1</intersection>
<intersection>-184.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-188,48.5,-188</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>48.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-184.5,53,-184.5</points>
<connection>
<GID>86</GID>
<name>IN_2</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-182.5,53,-182.5</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<connection>
<GID>86</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-180.5,48.5,-176</points>
<intersection>-180.5 2</intersection>
<intersection>-176 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-176,48.5,-176</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>48.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-180.5,53,-180.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,3.8147e-007,81.6,-91.8</PageViewport></page 1>
<page 2>
<PageViewport>0,3.8147e-007,81.6,-91.8</PageViewport></page 2>
<page 3>
<PageViewport>0,3.8147e-007,81.6,-91.8</PageViewport></page 3>
<page 4>
<PageViewport>0,3.8147e-007,81.6,-91.8</PageViewport></page 4>
<page 5>
<PageViewport>0,3.8147e-007,81.6,-91.8</PageViewport></page 5>
<page 6>
<PageViewport>0,3.8147e-007,81.6,-91.8</PageViewport></page 6>
<page 7>
<PageViewport>0,3.8147e-007,81.6,-91.8</PageViewport></page 7>
<page 8>
<PageViewport>0,3.8147e-007,81.6,-91.8</PageViewport></page 8>
<page 9>
<PageViewport>0,3.8147e-007,81.6,-91.8</PageViewport></page 9></circuit>