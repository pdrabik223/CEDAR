<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-105.285,-68.1114,111.325,-175.178</PageViewport>
<gate>
<ID>1</ID>
<type>AM_REGISTER16</type>
<position>8,-24</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>61 </input>
<input>
<ID>IN_10</ID>70 </input>
<input>
<ID>IN_11</ID>71 </input>
<input>
<ID>IN_12</ID>72 </input>
<input>
<ID>IN_13</ID>73 </input>
<input>
<ID>IN_14</ID>74 </input>
<input>
<ID>IN_15</ID>75 </input>
<input>
<ID>IN_2</ID>62 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_4</ID>64 </input>
<input>
<ID>IN_5</ID>65 </input>
<input>
<ID>IN_6</ID>66 </input>
<input>
<ID>IN_7</ID>67 </input>
<input>
<ID>IN_8</ID>68 </input>
<input>
<ID>IN_9</ID>69 </input>
<output>
<ID>OUT_0</ID>18 </output>
<output>
<ID>OUT_1</ID>13 </output>
<output>
<ID>OUT_10</ID>1 </output>
<output>
<ID>OUT_11</ID>12 </output>
<output>
<ID>OUT_12</ID>10 </output>
<output>
<ID>OUT_13</ID>16 </output>
<output>
<ID>OUT_14</ID>17 </output>
<output>
<ID>OUT_15</ID>3 </output>
<output>
<ID>OUT_2</ID>14 </output>
<output>
<ID>OUT_3</ID>7 </output>
<output>
<ID>OUT_4</ID>15 </output>
<output>
<ID>OUT_5</ID>8 </output>
<output>
<ID>OUT_6</ID>2 </output>
<output>
<ID>OUT_7</ID>19 </output>
<output>
<ID>OUT_8</ID>11 </output>
<output>
<ID>OUT_9</ID>9 </output>
<input>
<ID>clear</ID>82 </input>
<input>
<ID>clock</ID>77 </input>
<input>
<ID>load</ID>93 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 233</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>195</ID>
<type>AE_SMALL_INVERTER</type>
<position>-102,-78.5</position>
<input>
<ID>IN_0</ID>305 </input>
<output>
<ID>OUT_0</ID>304 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>126,-64.5</position>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_SMALL_INVERTER</type>
<position>7.5,-7</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>197</ID>
<type>AE_SMALL_INVERTER</type>
<position>-98,-78.5</position>
<input>
<ID>IN_0</ID>304 </input>
<output>
<ID>OUT_0</ID>309 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>113.5,-64.5</position>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>5</ID>
<type>BB_CLOCK</type>
<position>-124,-104</position>
<output>
<ID>CLK</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>17.5,-94.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>201</ID>
<type>BB_CLOCK</type>
<position>-114,-82.5</position>
<output>
<ID>CLK</ID>305 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_SMALL_INVERTER</type>
<position>7.5,-3</position>
<input>
<ID>IN_0</ID>23 </input>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_SMALL_INVERTER</type>
<position>7.5,1</position>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>203</ID>
<type>DA_FROM</type>
<position>-126,-77</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>10</ID>
<type>BB_CLOCK</type>
<position>-27.5,6</position>
<output>
<ID>CLK</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 25</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_SMALL_INVERTER</type>
<position>7.5,5</position>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>205</ID>
<type>DE_TO</type>
<position>-115,-98</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TO</lparam></gate>
<gate>
<ID>12</ID>
<type>AM_REGISTER16</type>
<position>18,-24</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_10</ID>1 </input>
<input>
<ID>IN_11</ID>12 </input>
<input>
<ID>IN_12</ID>10 </input>
<input>
<ID>IN_13</ID>16 </input>
<input>
<ID>IN_14</ID>17 </input>
<input>
<ID>IN_15</ID>3 </input>
<input>
<ID>IN_2</ID>14 </input>
<input>
<ID>IN_3</ID>7 </input>
<input>
<ID>IN_4</ID>15 </input>
<input>
<ID>IN_5</ID>8 </input>
<input>
<ID>IN_6</ID>2 </input>
<input>
<ID>IN_7</ID>19 </input>
<input>
<ID>IN_8</ID>11 </input>
<input>
<ID>IN_9</ID>9 </input>
<output>
<ID>OUT_0</ID>42 </output>
<output>
<ID>OUT_1</ID>43 </output>
<output>
<ID>OUT_10</ID>52 </output>
<output>
<ID>OUT_11</ID>53 </output>
<output>
<ID>OUT_12</ID>54 </output>
<output>
<ID>OUT_13</ID>55 </output>
<output>
<ID>OUT_14</ID>56 </output>
<output>
<ID>OUT_15</ID>57 </output>
<output>
<ID>OUT_2</ID>44 </output>
<output>
<ID>OUT_3</ID>45 </output>
<output>
<ID>OUT_4</ID>46 </output>
<output>
<ID>OUT_5</ID>47 </output>
<output>
<ID>OUT_6</ID>48 </output>
<output>
<ID>OUT_7</ID>49 </output>
<output>
<ID>OUT_8</ID>50 </output>
<output>
<ID>OUT_9</ID>51 </output>
<input>
<ID>clear</ID>82 </input>
<input>
<ID>clock</ID>101 </input>
<input>
<ID>count_enable</ID>98 </input>
<input>
<ID>load</ID>110 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 233</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>206</ID>
<type>DE_TO</type>
<position>-64,-78.5</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_OR2</type>
<position>7,-36.5</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>DE_TO</type>
<position>-90.5,-87.5</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2</lparam></gate>
<gate>
<ID>208</ID>
<type>AE_SMALL_INVERTER</type>
<position>-94,-78.5</position>
<input>
<ID>IN_0</ID>309 </input>
<output>
<ID>OUT_0</ID>314 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>-10.5,5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ck</lparam></gate>
<gate>
<ID>17</ID>
<type>DA_FROM</type>
<position>-13,-7.5</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ck</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>-1.5,5.5</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ck</lparam></gate>
<gate>
<ID>212</ID>
<type>AE_SMALL_INVERTER</type>
<position>-90,-78.5</position>
<input>
<ID>IN_0</ID>314 </input>
<output>
<ID>OUT_0</ID>316 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>4,-43.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ck</lparam></gate>
<gate>
<ID>213</ID>
<type>AE_SMALL_INVERTER</type>
<position>-86,-78.5</position>
<input>
<ID>IN_0</ID>316 </input>
<output>
<ID>OUT_0</ID>317 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_SMALL_INVERTER</type>
<position>-90,-106</position>
<input>
<ID>IN_0</ID>92 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>0,-14.5</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ck</lparam></gate>
<gate>
<ID>215</ID>
<type>AE_SMALL_INVERTER</type>
<position>-82,-78.5</position>
<input>
<ID>IN_0</ID>317 </input>
<output>
<ID>OUT_0</ID>318 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_SMALL_INVERTER</type>
<position>19.5,-8.5</position>
<input>
<ID>IN_0</ID>109 </input>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_FULLADDER_4BIT</type>
<position>58.5,-43</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>39 </input>
<input>
<ID>IN_3</ID>40 </input>
<input>
<ID>IN_B_0</ID>54 </input>
<input>
<ID>IN_B_1</ID>55 </input>
<input>
<ID>IN_B_2</ID>56 </input>
<input>
<ID>IN_B_3</ID>57 </input>
<output>
<ID>OUT_0</ID>72 </output>
<output>
<ID>OUT_1</ID>73 </output>
<output>
<ID>OUT_2</ID>74 </output>
<output>
<ID>OUT_3</ID>75 </output>
<input>
<ID>carry_in</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_FULLADDER_4BIT</type>
<position>74.5,-43</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>35 </input>
<input>
<ID>IN_3</ID>36 </input>
<input>
<ID>IN_B_0</ID>50 </input>
<input>
<ID>IN_B_1</ID>51 </input>
<input>
<ID>IN_B_2</ID>52 </input>
<input>
<ID>IN_B_3</ID>53 </input>
<output>
<ID>OUT_0</ID>68 </output>
<output>
<ID>OUT_1</ID>69 </output>
<output>
<ID>OUT_2</ID>70 </output>
<output>
<ID>OUT_3</ID>71 </output>
<input>
<ID>carry_in</ID>5 </input>
<output>
<ID>carry_out</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_FULLADDER_4BIT</type>
<position>90.5,-43</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>31 </input>
<input>
<ID>IN_3</ID>32 </input>
<input>
<ID>IN_B_0</ID>46 </input>
<input>
<ID>IN_B_1</ID>47 </input>
<input>
<ID>IN_B_2</ID>48 </input>
<input>
<ID>IN_B_3</ID>49 </input>
<output>
<ID>OUT_0</ID>64 </output>
<output>
<ID>OUT_1</ID>65 </output>
<output>
<ID>OUT_2</ID>66 </output>
<output>
<ID>OUT_3</ID>67 </output>
<input>
<ID>carry_in</ID>6 </input>
<output>
<ID>carry_out</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_FULLADDER_4BIT</type>
<position>106.5,-43</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<input>
<ID>IN_2</ID>27 </input>
<input>
<ID>IN_3</ID>28 </input>
<input>
<ID>IN_B_0</ID>42 </input>
<input>
<ID>IN_B_1</ID>43 </input>
<input>
<ID>IN_B_2</ID>44 </input>
<input>
<ID>IN_B_3</ID>45 </input>
<output>
<ID>OUT_0</ID>60 </output>
<output>
<ID>OUT_1</ID>61 </output>
<output>
<ID>OUT_2</ID>62 </output>
<output>
<ID>OUT_3</ID>63 </output>
<output>
<ID>carry_out</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>27</ID>
<type>AM_REGISTER16</type>
<position>42,-1.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_10</ID>52 </input>
<input>
<ID>IN_11</ID>53 </input>
<input>
<ID>IN_12</ID>54 </input>
<input>
<ID>IN_13</ID>55 </input>
<input>
<ID>IN_14</ID>56 </input>
<input>
<ID>IN_15</ID>57 </input>
<input>
<ID>IN_2</ID>44 </input>
<input>
<ID>IN_3</ID>45 </input>
<input>
<ID>IN_4</ID>46 </input>
<input>
<ID>IN_5</ID>47 </input>
<input>
<ID>IN_6</ID>48 </input>
<input>
<ID>IN_7</ID>49 </input>
<input>
<ID>IN_8</ID>50 </input>
<input>
<ID>IN_9</ID>51 </input>
<output>
<ID>OUT_0</ID>25 </output>
<output>
<ID>OUT_1</ID>26 </output>
<output>
<ID>OUT_10</ID>35 </output>
<output>
<ID>OUT_11</ID>36 </output>
<output>
<ID>OUT_12</ID>37 </output>
<output>
<ID>OUT_13</ID>38 </output>
<output>
<ID>OUT_14</ID>39 </output>
<output>
<ID>OUT_15</ID>40 </output>
<output>
<ID>OUT_2</ID>27 </output>
<output>
<ID>OUT_3</ID>28 </output>
<output>
<ID>OUT_4</ID>29 </output>
<output>
<ID>OUT_5</ID>30 </output>
<output>
<ID>OUT_6</ID>31 </output>
<output>
<ID>OUT_7</ID>32 </output>
<output>
<ID>OUT_8</ID>33 </output>
<output>
<ID>OUT_9</ID>34 </output>
<input>
<ID>clear</ID>82 </input>
<input>
<ID>clock</ID>100 </input>
<input>
<ID>load</ID>97 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 144</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_SMALL_INVERTER</type>
<position>19.5,-4.5</position>
<input>
<ID>IN_0</ID>99 </input>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>29</ID>
<type>CC_PULSE</type>
<position>-39.5,-11</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AE_SMALL_INVERTER</type>
<position>19.5,-0.5</position>
<input>
<ID>IN_0</ID>102 </input>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_REGISTER8</type>
<position>-1.5,-2.5</position>
<input>
<ID>clear</ID>82 </input>
<input>
<ID>clock</ID>79 </input>
<input>
<ID>count_enable</ID>87 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 12</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>32</ID>
<type>AE_SMALL_INVERTER</type>
<position>19.5,3.5</position>
<input>
<ID>IN_0</ID>103 </input>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>-19.5,-4</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_SMALL_INVERTER</type>
<position>22.5,5.5</position>
<input>
<ID>IN_0</ID>97 </input>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>-15.5,5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AE_SMALL_INVERTER</type>
<position>22.5,1.5</position>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>37</ID>
<type>AE_OR2</type>
<position>-8,-8.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AE_SMALL_INVERTER</type>
<position>22.5,-2.5</position>
<input>
<ID>IN_0</ID>106 </input>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>-19.5,6</position>
<input>
<ID>N_in0</ID>81 </input>
<input>
<ID>N_in1</ID>80 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AE_SMALL_INVERTER</type>
<position>22.5,-6.5</position>
<input>
<ID>IN_0</ID>105 </input>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>43</ID>
<type>AE_SMALL_INVERTER</type>
<position>10.5,7</position>
<input>
<ID>IN_0</ID>96 </input>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>44</ID>
<type>AE_SMALL_INVERTER</type>
<position>10.5,3</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_SMALL_INVERTER</type>
<position>10.5,-1</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>46</ID>
<type>AE_SMALL_INVERTER</type>
<position>10.5,-5</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_SMALL_INVERTER</type>
<position>-94,-106</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>52</ID>
<type>AM_RAM_16x16</type>
<position>3.5,-92.5</position>
<input>
<ID>ADDRESS_0</ID>115 </input>
<input>
<ID>ADDRESS_1</ID>116 </input>
<input>
<ID>ADDRESS_10</ID>123 </input>
<input>
<ID>ADDRESS_11</ID>124 </input>
<input>
<ID>ADDRESS_12</ID>125 </input>
<input>
<ID>ADDRESS_13</ID>119 </input>
<input>
<ID>ADDRESS_14</ID>120 </input>
<input>
<ID>ADDRESS_15</ID>121 </input>
<input>
<ID>ADDRESS_2</ID>117 </input>
<input>
<ID>ADDRESS_3</ID>113 </input>
<input>
<ID>ADDRESS_4</ID>112 </input>
<input>
<ID>ADDRESS_5</ID>114 </input>
<input>
<ID>ADDRESS_6</ID>118 </input>
<input>
<ID>ADDRESS_7</ID>127 </input>
<input>
<ID>ADDRESS_8</ID>126 </input>
<input>
<ID>ADDRESS_9</ID>122 </input>
<input>
<ID>DATA_IN_0</ID>179 </input>
<input>
<ID>DATA_IN_1</ID>180 </input>
<input>
<ID>DATA_IN_10</ID>189 </input>
<input>
<ID>DATA_IN_11</ID>190 </input>
<input>
<ID>DATA_IN_12</ID>194 </input>
<input>
<ID>DATA_IN_13</ID>193 </input>
<input>
<ID>DATA_IN_14</ID>192 </input>
<input>
<ID>DATA_IN_15</ID>191 </input>
<input>
<ID>DATA_IN_2</ID>181 </input>
<input>
<ID>DATA_IN_3</ID>182 </input>
<input>
<ID>DATA_IN_4</ID>183 </input>
<input>
<ID>DATA_IN_5</ID>184 </input>
<input>
<ID>DATA_IN_6</ID>185 </input>
<input>
<ID>DATA_IN_7</ID>186 </input>
<input>
<ID>DATA_IN_8</ID>187 </input>
<input>
<ID>DATA_IN_9</ID>188 </input>
<output>
<ID>DATA_OUT_0</ID>179 </output>
<output>
<ID>DATA_OUT_1</ID>180 </output>
<output>
<ID>DATA_OUT_10</ID>189 </output>
<output>
<ID>DATA_OUT_11</ID>190 </output>
<output>
<ID>DATA_OUT_12</ID>194 </output>
<output>
<ID>DATA_OUT_13</ID>193 </output>
<output>
<ID>DATA_OUT_14</ID>192 </output>
<output>
<ID>DATA_OUT_15</ID>191 </output>
<output>
<ID>DATA_OUT_2</ID>181 </output>
<output>
<ID>DATA_OUT_3</ID>182 </output>
<output>
<ID>DATA_OUT_4</ID>183 </output>
<output>
<ID>DATA_OUT_5</ID>184 </output>
<output>
<ID>DATA_OUT_6</ID>185 </output>
<output>
<ID>DATA_OUT_7</ID>186 </output>
<output>
<ID>DATA_OUT_8</ID>187 </output>
<output>
<ID>DATA_OUT_9</ID>188 </output>
<input>
<ID>write_clock</ID>134 </input>
<input>
<ID>write_enable</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 16</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:1 1</lparam>
<lparam>Address:2 2</lparam>
<lparam>Address:3 3</lparam>
<lparam>Address:4 4</lparam>
<lparam>Address:5 5</lparam>
<lparam>Address:6 6</lparam>
<lparam>Address:7 7</lparam>
<lparam>Address:8 8</lparam>
<lparam>Address:9 9</lparam>
<lparam>Address:10 16</lparam>
<lparam>Address:11 17</lparam>
<lparam>Address:12 18</lparam>
<lparam>Address:13 19</lparam>
<lparam>Address:14 20</lparam>
<lparam>Address:15 21</lparam>
<lparam>Address:16 22</lparam>
<lparam>Address:17 23</lparam>
<lparam>Address:18 24</lparam>
<lparam>Address:19 25</lparam>
<lparam>Address:20 32</lparam>
<lparam>Address:21 33</lparam>
<lparam>Address:22 34</lparam>
<lparam>Address:23 35</lparam>
<lparam>Address:24 36</lparam>
<lparam>Address:25 37</lparam>
<lparam>Address:26 38</lparam>
<lparam>Address:27 39</lparam>
<lparam>Address:28 40</lparam>
<lparam>Address:29 41</lparam>
<lparam>Address:30 48</lparam>
<lparam>Address:31 49</lparam>
<lparam>Address:32 50</lparam>
<lparam>Address:33 51</lparam>
<lparam>Address:34 52</lparam>
<lparam>Address:35 53</lparam>
<lparam>Address:36 54</lparam>
<lparam>Address:37 55</lparam>
<lparam>Address:38 56</lparam>
<lparam>Address:39 57</lparam>
<lparam>Address:40 64</lparam>
<lparam>Address:41 65</lparam>
<lparam>Address:42 66</lparam>
<lparam>Address:43 67</lparam>
<lparam>Address:44 68</lparam>
<lparam>Address:45 69</lparam>
<lparam>Address:46 70</lparam>
<lparam>Address:47 71</lparam>
<lparam>Address:48 72</lparam>
<lparam>Address:49 73</lparam>
<lparam>Address:50 80</lparam>
<lparam>Address:51 81</lparam>
<lparam>Address:52 82</lparam>
<lparam>Address:53 83</lparam>
<lparam>Address:54 84</lparam>
<lparam>Address:55 85</lparam>
<lparam>Address:56 86</lparam>
<lparam>Address:57 87</lparam>
<lparam>Address:58 88</lparam>
<lparam>Address:59 89</lparam>
<lparam>Address:60 96</lparam>
<lparam>Address:61 97</lparam>
<lparam>Address:62 98</lparam>
<lparam>Address:63 99</lparam>
<lparam>Address:64 100</lparam>
<lparam>Address:65 101</lparam>
<lparam>Address:66 102</lparam>
<lparam>Address:67 103</lparam>
<lparam>Address:68 104</lparam>
<lparam>Address:69 105</lparam>
<lparam>Address:70 112</lparam>
<lparam>Address:71 113</lparam>
<lparam>Address:72 114</lparam>
<lparam>Address:73 115</lparam>
<lparam>Address:74 116</lparam>
<lparam>Address:75 117</lparam>
<lparam>Address:76 118</lparam>
<lparam>Address:77 119</lparam>
<lparam>Address:78 120</lparam>
<lparam>Address:79 121</lparam>
<lparam>Address:80 128</lparam>
<lparam>Address:81 129</lparam>
<lparam>Address:82 130</lparam>
<lparam>Address:83 131</lparam>
<lparam>Address:84 132</lparam>
<lparam>Address:85 133</lparam>
<lparam>Address:86 134</lparam>
<lparam>Address:87 135</lparam>
<lparam>Address:88 136</lparam>
<lparam>Address:89 137</lparam>
<lparam>Address:90 144</lparam>
<lparam>Address:91 145</lparam>
<lparam>Address:92 146</lparam>
<lparam>Address:93 147</lparam>
<lparam>Address:94 148</lparam>
<lparam>Address:95 149</lparam>
<lparam>Address:96 150</lparam>
<lparam>Address:97 151</lparam>
<lparam>Address:98 152</lparam>
<lparam>Address:99 153</lparam>
<lparam>Address:100 256</lparam>
<lparam>Address:101 257</lparam>
<lparam>Address:102 258</lparam>
<lparam>Address:103 259</lparam>
<lparam>Address:104 260</lparam>
<lparam>Address:105 261</lparam>
<lparam>Address:106 262</lparam>
<lparam>Address:107 263</lparam>
<lparam>Address:108 264</lparam>
<lparam>Address:109 265</lparam>
<lparam>Address:110 272</lparam>
<lparam>Address:111 273</lparam>
<lparam>Address:112 274</lparam>
<lparam>Address:113 275</lparam>
<lparam>Address:114 276</lparam>
<lparam>Address:115 277</lparam>
<lparam>Address:116 278</lparam>
<lparam>Address:117 279</lparam>
<lparam>Address:118 280</lparam>
<lparam>Address:119 281</lparam>
<lparam>Address:120 288</lparam>
<lparam>Address:121 289</lparam>
<lparam>Address:122 290</lparam>
<lparam>Address:123 291</lparam>
<lparam>Address:124 292</lparam>
<lparam>Address:125 293</lparam>
<lparam>Address:126 294</lparam>
<lparam>Address:127 295</lparam>
<lparam>Address:128 296</lparam>
<lparam>Address:129 297</lparam>
<lparam>Address:130 304</lparam>
<lparam>Address:131 305</lparam>
<lparam>Address:132 306</lparam>
<lparam>Address:133 307</lparam>
<lparam>Address:134 308</lparam>
<lparam>Address:135 309</lparam>
<lparam>Address:136 310</lparam>
<lparam>Address:137 311</lparam>
<lparam>Address:138 312</lparam>
<lparam>Address:139 313</lparam>
<lparam>Address:140 320</lparam>
<lparam>Address:141 321</lparam>
<lparam>Address:142 322</lparam>
<lparam>Address:143 323</lparam>
<lparam>Address:144 324</lparam>
<lparam>Address:145 325</lparam>
<lparam>Address:146 326</lparam>
<lparam>Address:147 327</lparam>
<lparam>Address:148 328</lparam>
<lparam>Address:149 329</lparam>
<lparam>Address:150 336</lparam>
<lparam>Address:151 337</lparam>
<lparam>Address:152 338</lparam>
<lparam>Address:153 339</lparam>
<lparam>Address:154 340</lparam>
<lparam>Address:155 341</lparam>
<lparam>Address:156 342</lparam>
<lparam>Address:157 343</lparam>
<lparam>Address:158 344</lparam>
<lparam>Address:159 345</lparam>
<lparam>Address:160 352</lparam>
<lparam>Address:161 353</lparam>
<lparam>Address:162 354</lparam>
<lparam>Address:163 355</lparam>
<lparam>Address:164 356</lparam>
<lparam>Address:165 357</lparam>
<lparam>Address:166 358</lparam>
<lparam>Address:167 359</lparam>
<lparam>Address:168 360</lparam>
<lparam>Address:169 361</lparam>
<lparam>Address:170 368</lparam>
<lparam>Address:171 369</lparam>
<lparam>Address:172 370</lparam>
<lparam>Address:173 371</lparam>
<lparam>Address:174 372</lparam>
<lparam>Address:175 373</lparam>
<lparam>Address:176 374</lparam>
<lparam>Address:177 375</lparam>
<lparam>Address:178 376</lparam>
<lparam>Address:179 377</lparam>
<lparam>Address:180 384</lparam>
<lparam>Address:181 385</lparam>
<lparam>Address:182 386</lparam>
<lparam>Address:183 387</lparam>
<lparam>Address:184 388</lparam>
<lparam>Address:185 389</lparam>
<lparam>Address:186 390</lparam>
<lparam>Address:187 391</lparam>
<lparam>Address:188 392</lparam>
<lparam>Address:189 393</lparam>
<lparam>Address:190 400</lparam>
<lparam>Address:191 401</lparam>
<lparam>Address:192 402</lparam>
<lparam>Address:193 403</lparam>
<lparam>Address:194 404</lparam>
<lparam>Address:195 405</lparam>
<lparam>Address:196 406</lparam>
<lparam>Address:197 407</lparam>
<lparam>Address:198 408</lparam>
<lparam>Address:199 409</lparam>
<lparam>Address:200 512</lparam>
<lparam>Address:201 513</lparam>
<lparam>Address:202 514</lparam>
<lparam>Address:203 515</lparam>
<lparam>Address:204 516</lparam>
<lparam>Address:205 517</lparam>
<lparam>Address:206 518</lparam>
<lparam>Address:207 519</lparam>
<lparam>Address:208 520</lparam>
<lparam>Address:209 521</lparam>
<lparam>Address:210 528</lparam>
<lparam>Address:211 529</lparam>
<lparam>Address:212 530</lparam>
<lparam>Address:213 531</lparam>
<lparam>Address:214 532</lparam>
<lparam>Address:215 533</lparam>
<lparam>Address:216 534</lparam>
<lparam>Address:217 535</lparam>
<lparam>Address:218 536</lparam>
<lparam>Address:219 537</lparam>
<lparam>Address:220 544</lparam>
<lparam>Address:221 545</lparam>
<lparam>Address:222 546</lparam>
<lparam>Address:223 547</lparam>
<lparam>Address:224 548</lparam>
<lparam>Address:225 549</lparam>
<lparam>Address:226 550</lparam>
<lparam>Address:227 551</lparam>
<lparam>Address:228 552</lparam>
<lparam>Address:229 553</lparam>
<lparam>Address:230 560</lparam>
<lparam>Address:231 561</lparam>
<lparam>Address:232 562</lparam>
<lparam>Address:233 563</lparam>
<lparam>Address:234 564</lparam>
<lparam>Address:235 565</lparam>
<lparam>Address:236 566</lparam>
<lparam>Address:237 567</lparam>
<lparam>Address:238 568</lparam>
<lparam>Address:239 569</lparam>
<lparam>Address:240 576</lparam>
<lparam>Address:241 577</lparam>
<lparam>Address:242 578</lparam>
<lparam>Address:243 579</lparam>
<lparam>Address:244 580</lparam>
<lparam>Address:245 581</lparam>
<lparam>Address:246 582</lparam>
<lparam>Address:247 583</lparam>
<lparam>Address:248 584</lparam>
<lparam>Address:249 585</lparam>
<lparam>Address:250 592</lparam>
<lparam>Address:251 593</lparam>
<lparam>Address:252 594</lparam>
<lparam>Address:253 595</lparam>
<lparam>Address:254 596</lparam>
<lparam>Address:255 597</lparam>
<lparam>Address:256 598</lparam>
<lparam>Address:257 599</lparam>
<lparam>Address:258 600</lparam>
<lparam>Address:259 601</lparam>
<lparam>Address:260 608</lparam>
<lparam>Address:261 609</lparam>
<lparam>Address:262 610</lparam>
<lparam>Address:263 611</lparam>
<lparam>Address:264 612</lparam>
<lparam>Address:265 613</lparam>
<lparam>Address:266 614</lparam>
<lparam>Address:267 615</lparam>
<lparam>Address:268 616</lparam>
<lparam>Address:269 617</lparam>
<lparam>Address:270 624</lparam>
<lparam>Address:271 625</lparam>
<lparam>Address:272 626</lparam>
<lparam>Address:273 627</lparam>
<lparam>Address:274 628</lparam>
<lparam>Address:275 629</lparam>
<lparam>Address:276 630</lparam>
<lparam>Address:277 631</lparam>
<lparam>Address:278 632</lparam>
<lparam>Address:279 633</lparam>
<lparam>Address:280 640</lparam>
<lparam>Address:281 641</lparam>
<lparam>Address:282 642</lparam>
<lparam>Address:283 643</lparam>
<lparam>Address:284 644</lparam>
<lparam>Address:285 645</lparam>
<lparam>Address:286 646</lparam>
<lparam>Address:287 647</lparam>
<lparam>Address:288 648</lparam>
<lparam>Address:289 649</lparam>
<lparam>Address:290 656</lparam>
<lparam>Address:291 657</lparam>
<lparam>Address:292 658</lparam>
<lparam>Address:293 659</lparam>
<lparam>Address:294 660</lparam>
<lparam>Address:295 661</lparam>
<lparam>Address:296 662</lparam>
<lparam>Address:297 663</lparam>
<lparam>Address:298 664</lparam>
<lparam>Address:299 665</lparam>
<lparam>Address:300 768</lparam>
<lparam>Address:301 769</lparam>
<lparam>Address:302 770</lparam>
<lparam>Address:303 771</lparam>
<lparam>Address:304 772</lparam>
<lparam>Address:305 773</lparam>
<lparam>Address:306 774</lparam>
<lparam>Address:307 775</lparam>
<lparam>Address:308 776</lparam>
<lparam>Address:309 777</lparam>
<lparam>Address:310 784</lparam>
<lparam>Address:311 785</lparam>
<lparam>Address:312 786</lparam>
<lparam>Address:313 787</lparam>
<lparam>Address:314 788</lparam>
<lparam>Address:315 789</lparam>
<lparam>Address:316 790</lparam>
<lparam>Address:317 791</lparam>
<lparam>Address:318 792</lparam>
<lparam>Address:319 793</lparam>
<lparam>Address:320 800</lparam>
<lparam>Address:321 801</lparam>
<lparam>Address:322 802</lparam>
<lparam>Address:323 803</lparam>
<lparam>Address:324 804</lparam>
<lparam>Address:325 805</lparam>
<lparam>Address:326 806</lparam>
<lparam>Address:327 807</lparam>
<lparam>Address:328 808</lparam>
<lparam>Address:329 809</lparam>
<lparam>Address:330 816</lparam>
<lparam>Address:331 817</lparam>
<lparam>Address:332 818</lparam>
<lparam>Address:333 819</lparam>
<lparam>Address:334 820</lparam>
<lparam>Address:335 821</lparam>
<lparam>Address:336 822</lparam>
<lparam>Address:337 823</lparam>
<lparam>Address:338 824</lparam>
<lparam>Address:339 825</lparam>
<lparam>Address:340 832</lparam>
<lparam>Address:341 833</lparam>
<lparam>Address:342 834</lparam>
<lparam>Address:343 835</lparam>
<lparam>Address:344 836</lparam>
<lparam>Address:345 837</lparam>
<lparam>Address:346 838</lparam>
<lparam>Address:347 839</lparam>
<lparam>Address:348 840</lparam>
<lparam>Address:349 841</lparam>
<lparam>Address:350 848</lparam>
<lparam>Address:351 849</lparam>
<lparam>Address:352 850</lparam>
<lparam>Address:353 851</lparam>
<lparam>Address:354 852</lparam>
<lparam>Address:355 853</lparam>
<lparam>Address:356 854</lparam>
<lparam>Address:357 855</lparam>
<lparam>Address:358 856</lparam>
<lparam>Address:359 857</lparam>
<lparam>Address:360 864</lparam>
<lparam>Address:361 865</lparam>
<lparam>Address:362 866</lparam>
<lparam>Address:363 867</lparam>
<lparam>Address:364 868</lparam>
<lparam>Address:365 869</lparam>
<lparam>Address:366 870</lparam>
<lparam>Address:367 871</lparam>
<lparam>Address:368 872</lparam>
<lparam>Address:369 873</lparam>
<lparam>Address:370 880</lparam>
<lparam>Address:371 881</lparam>
<lparam>Address:372 882</lparam>
<lparam>Address:373 883</lparam>
<lparam>Address:374 884</lparam>
<lparam>Address:375 885</lparam>
<lparam>Address:376 886</lparam>
<lparam>Address:377 887</lparam>
<lparam>Address:378 888</lparam>
<lparam>Address:379 889</lparam>
<lparam>Address:380 896</lparam>
<lparam>Address:381 897</lparam>
<lparam>Address:382 898</lparam>
<lparam>Address:383 899</lparam>
<lparam>Address:384 900</lparam>
<lparam>Address:385 901</lparam>
<lparam>Address:386 902</lparam>
<lparam>Address:387 903</lparam>
<lparam>Address:388 904</lparam>
<lparam>Address:389 905</lparam>
<lparam>Address:390 912</lparam>
<lparam>Address:391 913</lparam>
<lparam>Address:392 914</lparam>
<lparam>Address:393 915</lparam>
<lparam>Address:394 916</lparam>
<lparam>Address:395 917</lparam>
<lparam>Address:396 918</lparam>
<lparam>Address:397 919</lparam>
<lparam>Address:398 920</lparam>
<lparam>Address:399 921</lparam>
<lparam>Address:400 1024</lparam>
<lparam>Address:401 1025</lparam>
<lparam>Address:402 1026</lparam>
<lparam>Address:403 1027</lparam>
<lparam>Address:404 1028</lparam>
<lparam>Address:405 1029</lparam>
<lparam>Address:406 1030</lparam>
<lparam>Address:407 1031</lparam>
<lparam>Address:408 1032</lparam>
<lparam>Address:409 1033</lparam>
<lparam>Address:410 1040</lparam>
<lparam>Address:411 1041</lparam>
<lparam>Address:412 1042</lparam>
<lparam>Address:413 1043</lparam>
<lparam>Address:414 1044</lparam>
<lparam>Address:415 1045</lparam>
<lparam>Address:416 1046</lparam>
<lparam>Address:417 1047</lparam>
<lparam>Address:418 1048</lparam>
<lparam>Address:419 1049</lparam>
<lparam>Address:420 1056</lparam>
<lparam>Address:421 1057</lparam>
<lparam>Address:422 1058</lparam>
<lparam>Address:423 1059</lparam>
<lparam>Address:424 1060</lparam>
<lparam>Address:425 1061</lparam>
<lparam>Address:426 1062</lparam>
<lparam>Address:427 1063</lparam>
<lparam>Address:428 1064</lparam>
<lparam>Address:429 1065</lparam>
<lparam>Address:430 1072</lparam>
<lparam>Address:431 1073</lparam>
<lparam>Address:432 1074</lparam>
<lparam>Address:433 1075</lparam>
<lparam>Address:434 1076</lparam>
<lparam>Address:435 1077</lparam>
<lparam>Address:436 1078</lparam>
<lparam>Address:437 1079</lparam>
<lparam>Address:438 1080</lparam>
<lparam>Address:439 1081</lparam>
<lparam>Address:440 1088</lparam>
<lparam>Address:441 1089</lparam>
<lparam>Address:442 1090</lparam>
<lparam>Address:443 1091</lparam>
<lparam>Address:444 1092</lparam>
<lparam>Address:445 1093</lparam>
<lparam>Address:446 1094</lparam>
<lparam>Address:447 1095</lparam>
<lparam>Address:448 1096</lparam>
<lparam>Address:449 1097</lparam>
<lparam>Address:450 1104</lparam>
<lparam>Address:451 1105</lparam>
<lparam>Address:452 1106</lparam>
<lparam>Address:453 1107</lparam>
<lparam>Address:454 1108</lparam>
<lparam>Address:455 1109</lparam>
<lparam>Address:456 1110</lparam>
<lparam>Address:457 1111</lparam>
<lparam>Address:458 1112</lparam>
<lparam>Address:459 1113</lparam>
<lparam>Address:460 1120</lparam>
<lparam>Address:461 1121</lparam>
<lparam>Address:462 1122</lparam>
<lparam>Address:463 1123</lparam>
<lparam>Address:464 1124</lparam>
<lparam>Address:465 1125</lparam>
<lparam>Address:466 1126</lparam>
<lparam>Address:467 1127</lparam>
<lparam>Address:468 1128</lparam>
<lparam>Address:469 1129</lparam>
<lparam>Address:470 1136</lparam>
<lparam>Address:471 1137</lparam>
<lparam>Address:472 1138</lparam>
<lparam>Address:473 1139</lparam>
<lparam>Address:474 1140</lparam>
<lparam>Address:475 1141</lparam>
<lparam>Address:476 1142</lparam>
<lparam>Address:477 1143</lparam>
<lparam>Address:478 1144</lparam>
<lparam>Address:479 1145</lparam>
<lparam>Address:480 1152</lparam>
<lparam>Address:481 1153</lparam>
<lparam>Address:482 1154</lparam>
<lparam>Address:483 1155</lparam>
<lparam>Address:484 1156</lparam>
<lparam>Address:485 1157</lparam>
<lparam>Address:486 1158</lparam>
<lparam>Address:487 1159</lparam>
<lparam>Address:488 1160</lparam>
<lparam>Address:489 1161</lparam>
<lparam>Address:490 1168</lparam>
<lparam>Address:491 1169</lparam>
<lparam>Address:492 1170</lparam>
<lparam>Address:493 1171</lparam>
<lparam>Address:494 1172</lparam>
<lparam>Address:495 1173</lparam>
<lparam>Address:496 1174</lparam>
<lparam>Address:497 1175</lparam>
<lparam>Address:498 1176</lparam>
<lparam>Address:499 1177</lparam>
<lparam>Address:500 1280</lparam>
<lparam>Address:501 1281</lparam>
<lparam>Address:502 1282</lparam>
<lparam>Address:503 1283</lparam>
<lparam>Address:504 1284</lparam>
<lparam>Address:505 1285</lparam>
<lparam>Address:506 1286</lparam>
<lparam>Address:507 1287</lparam>
<lparam>Address:508 1288</lparam>
<lparam>Address:509 1289</lparam>
<lparam>Address:510 1296</lparam>
<lparam>Address:511 1297</lparam>
<lparam>Address:512 1298</lparam>
<lparam>Address:513 1299</lparam>
<lparam>Address:514 1300</lparam>
<lparam>Address:515 1301</lparam>
<lparam>Address:516 1302</lparam>
<lparam>Address:517 1303</lparam>
<lparam>Address:518 1304</lparam>
<lparam>Address:519 1305</lparam>
<lparam>Address:520 1312</lparam>
<lparam>Address:521 1313</lparam>
<lparam>Address:522 1314</lparam>
<lparam>Address:523 1315</lparam>
<lparam>Address:524 1316</lparam>
<lparam>Address:525 1317</lparam>
<lparam>Address:526 1318</lparam>
<lparam>Address:527 1319</lparam>
<lparam>Address:528 1320</lparam>
<lparam>Address:529 1321</lparam>
<lparam>Address:530 1328</lparam>
<lparam>Address:531 1329</lparam>
<lparam>Address:532 1330</lparam>
<lparam>Address:533 1331</lparam>
<lparam>Address:534 1332</lparam>
<lparam>Address:535 1333</lparam>
<lparam>Address:536 1334</lparam>
<lparam>Address:537 1335</lparam>
<lparam>Address:538 1336</lparam>
<lparam>Address:539 1337</lparam>
<lparam>Address:540 1344</lparam>
<lparam>Address:541 1345</lparam>
<lparam>Address:542 1346</lparam>
<lparam>Address:543 1347</lparam>
<lparam>Address:544 1348</lparam>
<lparam>Address:545 1349</lparam>
<lparam>Address:546 1350</lparam>
<lparam>Address:547 1351</lparam>
<lparam>Address:548 1352</lparam>
<lparam>Address:549 1353</lparam>
<lparam>Address:550 1360</lparam>
<lparam>Address:551 1361</lparam>
<lparam>Address:552 1362</lparam>
<lparam>Address:553 1363</lparam>
<lparam>Address:554 1364</lparam>
<lparam>Address:555 1365</lparam>
<lparam>Address:556 1366</lparam>
<lparam>Address:557 1367</lparam>
<lparam>Address:558 1368</lparam>
<lparam>Address:559 1369</lparam>
<lparam>Address:560 1376</lparam>
<lparam>Address:561 1377</lparam>
<lparam>Address:562 1378</lparam>
<lparam>Address:563 1379</lparam>
<lparam>Address:564 1380</lparam>
<lparam>Address:565 1381</lparam>
<lparam>Address:566 1382</lparam>
<lparam>Address:567 1383</lparam>
<lparam>Address:568 1384</lparam>
<lparam>Address:569 1385</lparam>
<lparam>Address:570 1392</lparam>
<lparam>Address:571 1393</lparam>
<lparam>Address:572 1394</lparam>
<lparam>Address:573 1395</lparam>
<lparam>Address:574 1396</lparam>
<lparam>Address:575 1397</lparam>
<lparam>Address:576 1398</lparam>
<lparam>Address:577 1399</lparam>
<lparam>Address:578 1400</lparam>
<lparam>Address:579 1401</lparam>
<lparam>Address:580 1408</lparam>
<lparam>Address:581 1409</lparam>
<lparam>Address:582 1410</lparam>
<lparam>Address:583 1411</lparam>
<lparam>Address:584 1412</lparam>
<lparam>Address:585 1413</lparam>
<lparam>Address:586 1414</lparam>
<lparam>Address:587 1415</lparam>
<lparam>Address:588 1416</lparam>
<lparam>Address:589 1417</lparam>
<lparam>Address:590 1424</lparam>
<lparam>Address:591 1425</lparam>
<lparam>Address:592 1426</lparam>
<lparam>Address:593 1427</lparam>
<lparam>Address:594 1428</lparam>
<lparam>Address:595 1429</lparam>
<lparam>Address:596 1430</lparam>
<lparam>Address:597 1431</lparam>
<lparam>Address:598 1432</lparam>
<lparam>Address:599 1433</lparam>
<lparam>Address:600 1536</lparam>
<lparam>Address:601 1537</lparam>
<lparam>Address:602 1538</lparam>
<lparam>Address:603 1539</lparam>
<lparam>Address:604 1540</lparam>
<lparam>Address:605 1541</lparam>
<lparam>Address:606 1542</lparam>
<lparam>Address:607 1543</lparam>
<lparam>Address:608 1544</lparam>
<lparam>Address:609 1545</lparam>
<lparam>Address:610 1552</lparam>
<lparam>Address:611 1553</lparam>
<lparam>Address:612 1554</lparam>
<lparam>Address:613 1555</lparam>
<lparam>Address:614 1556</lparam>
<lparam>Address:615 1557</lparam>
<lparam>Address:616 1558</lparam>
<lparam>Address:617 1559</lparam>
<lparam>Address:618 1560</lparam>
<lparam>Address:619 1561</lparam>
<lparam>Address:620 1568</lparam>
<lparam>Address:621 1569</lparam>
<lparam>Address:622 1570</lparam>
<lparam>Address:623 1571</lparam>
<lparam>Address:624 1572</lparam>
<lparam>Address:625 1573</lparam>
<lparam>Address:626 1574</lparam>
<lparam>Address:627 1575</lparam>
<lparam>Address:628 1576</lparam>
<lparam>Address:629 1577</lparam>
<lparam>Address:630 1584</lparam>
<lparam>Address:631 1585</lparam>
<lparam>Address:632 1586</lparam>
<lparam>Address:633 1587</lparam>
<lparam>Address:634 1588</lparam>
<lparam>Address:635 1589</lparam>
<lparam>Address:636 1590</lparam>
<lparam>Address:637 1591</lparam>
<lparam>Address:638 1592</lparam>
<lparam>Address:639 1593</lparam>
<lparam>Address:640 1600</lparam>
<lparam>Address:641 1601</lparam>
<lparam>Address:642 1602</lparam>
<lparam>Address:643 1603</lparam>
<lparam>Address:644 1604</lparam>
<lparam>Address:645 1605</lparam>
<lparam>Address:646 1606</lparam>
<lparam>Address:647 1607</lparam>
<lparam>Address:648 1608</lparam>
<lparam>Address:649 1609</lparam>
<lparam>Address:650 1616</lparam>
<lparam>Address:651 1617</lparam>
<lparam>Address:652 1618</lparam>
<lparam>Address:653 1619</lparam>
<lparam>Address:654 1620</lparam>
<lparam>Address:655 1621</lparam>
<lparam>Address:656 1622</lparam>
<lparam>Address:657 1623</lparam>
<lparam>Address:658 1624</lparam>
<lparam>Address:659 1625</lparam>
<lparam>Address:660 1632</lparam>
<lparam>Address:661 1633</lparam>
<lparam>Address:662 1634</lparam>
<lparam>Address:663 1635</lparam>
<lparam>Address:664 1636</lparam>
<lparam>Address:665 1637</lparam>
<lparam>Address:666 1638</lparam>
<lparam>Address:667 1639</lparam>
<lparam>Address:668 1640</lparam>
<lparam>Address:669 1641</lparam>
<lparam>Address:670 1648</lparam>
<lparam>Address:671 1649</lparam>
<lparam>Address:672 1650</lparam>
<lparam>Address:673 1651</lparam>
<lparam>Address:674 1652</lparam>
<lparam>Address:675 1653</lparam>
<lparam>Address:676 1654</lparam>
<lparam>Address:677 1655</lparam>
<lparam>Address:678 1656</lparam>
<lparam>Address:679 1657</lparam>
<lparam>Address:680 1664</lparam>
<lparam>Address:681 1665</lparam>
<lparam>Address:682 1666</lparam>
<lparam>Address:683 1667</lparam>
<lparam>Address:684 1668</lparam>
<lparam>Address:685 1669</lparam>
<lparam>Address:686 1670</lparam>
<lparam>Address:687 1671</lparam>
<lparam>Address:688 1672</lparam>
<lparam>Address:689 1673</lparam>
<lparam>Address:690 1680</lparam>
<lparam>Address:691 1681</lparam>
<lparam>Address:692 1682</lparam>
<lparam>Address:693 1683</lparam>
<lparam>Address:694 1684</lparam>
<lparam>Address:695 1685</lparam>
<lparam>Address:696 1686</lparam>
<lparam>Address:697 1687</lparam>
<lparam>Address:698 1688</lparam>
<lparam>Address:699 1689</lparam>
<lparam>Address:700 1792</lparam>
<lparam>Address:701 1793</lparam>
<lparam>Address:702 1794</lparam>
<lparam>Address:703 1795</lparam>
<lparam>Address:704 1796</lparam>
<lparam>Address:705 1797</lparam>
<lparam>Address:706 1798</lparam>
<lparam>Address:707 1799</lparam>
<lparam>Address:708 1800</lparam>
<lparam>Address:709 1801</lparam>
<lparam>Address:710 1808</lparam>
<lparam>Address:711 1809</lparam>
<lparam>Address:712 1810</lparam>
<lparam>Address:713 1811</lparam>
<lparam>Address:714 1812</lparam>
<lparam>Address:715 1813</lparam>
<lparam>Address:716 1814</lparam>
<lparam>Address:717 1815</lparam>
<lparam>Address:718 1816</lparam>
<lparam>Address:719 1817</lparam>
<lparam>Address:720 1824</lparam>
<lparam>Address:721 1825</lparam>
<lparam>Address:722 1826</lparam>
<lparam>Address:723 1827</lparam>
<lparam>Address:724 1828</lparam>
<lparam>Address:725 1829</lparam>
<lparam>Address:726 1830</lparam>
<lparam>Address:727 1831</lparam>
<lparam>Address:728 1832</lparam>
<lparam>Address:729 1833</lparam>
<lparam>Address:730 1840</lparam>
<lparam>Address:731 1841</lparam>
<lparam>Address:732 1842</lparam>
<lparam>Address:733 1843</lparam>
<lparam>Address:734 1844</lparam>
<lparam>Address:735 1845</lparam>
<lparam>Address:736 1846</lparam>
<lparam>Address:737 1847</lparam>
<lparam>Address:738 1848</lparam>
<lparam>Address:739 1849</lparam>
<lparam>Address:740 1856</lparam>
<lparam>Address:741 1857</lparam>
<lparam>Address:742 1858</lparam>
<lparam>Address:743 1859</lparam>
<lparam>Address:744 1860</lparam>
<lparam>Address:745 1861</lparam>
<lparam>Address:746 1862</lparam>
<lparam>Address:747 1863</lparam>
<lparam>Address:748 1864</lparam>
<lparam>Address:749 1865</lparam>
<lparam>Address:750 1872</lparam>
<lparam>Address:751 1873</lparam>
<lparam>Address:752 1874</lparam>
<lparam>Address:753 1875</lparam>
<lparam>Address:754 1876</lparam>
<lparam>Address:755 1877</lparam>
<lparam>Address:756 1878</lparam>
<lparam>Address:757 1879</lparam>
<lparam>Address:758 1880</lparam>
<lparam>Address:759 1881</lparam>
<lparam>Address:760 1888</lparam>
<lparam>Address:761 1889</lparam>
<lparam>Address:762 1890</lparam>
<lparam>Address:763 1891</lparam>
<lparam>Address:764 1892</lparam>
<lparam>Address:765 1893</lparam>
<lparam>Address:766 1894</lparam>
<lparam>Address:767 1895</lparam>
<lparam>Address:768 1896</lparam>
<lparam>Address:769 1897</lparam>
<lparam>Address:770 1904</lparam>
<lparam>Address:771 1905</lparam>
<lparam>Address:772 1906</lparam>
<lparam>Address:773 1907</lparam>
<lparam>Address:774 1908</lparam>
<lparam>Address:775 1909</lparam>
<lparam>Address:776 1910</lparam>
<lparam>Address:777 1911</lparam>
<lparam>Address:778 1912</lparam>
<lparam>Address:779 1913</lparam>
<lparam>Address:780 1920</lparam>
<lparam>Address:781 1921</lparam>
<lparam>Address:782 1922</lparam>
<lparam>Address:783 1923</lparam>
<lparam>Address:784 1924</lparam>
<lparam>Address:785 1925</lparam>
<lparam>Address:786 1926</lparam>
<lparam>Address:787 1927</lparam>
<lparam>Address:788 1928</lparam>
<lparam>Address:789 1929</lparam>
<lparam>Address:790 1936</lparam>
<lparam>Address:791 1937</lparam>
<lparam>Address:792 1938</lparam>
<lparam>Address:793 1939</lparam>
<lparam>Address:794 1940</lparam>
<lparam>Address:795 1941</lparam>
<lparam>Address:796 1942</lparam>
<lparam>Address:797 1943</lparam>
<lparam>Address:798 1944</lparam>
<lparam>Address:799 1945</lparam>
<lparam>Address:800 2048</lparam>
<lparam>Address:801 2049</lparam>
<lparam>Address:802 2050</lparam>
<lparam>Address:803 2051</lparam>
<lparam>Address:804 2052</lparam>
<lparam>Address:805 2053</lparam>
<lparam>Address:806 2054</lparam>
<lparam>Address:807 2055</lparam>
<lparam>Address:808 2056</lparam>
<lparam>Address:809 2057</lparam>
<lparam>Address:810 2064</lparam>
<lparam>Address:811 2065</lparam>
<lparam>Address:812 2066</lparam>
<lparam>Address:813 2067</lparam>
<lparam>Address:814 2068</lparam>
<lparam>Address:815 2069</lparam>
<lparam>Address:816 2070</lparam>
<lparam>Address:817 2071</lparam>
<lparam>Address:818 2072</lparam>
<lparam>Address:819 2073</lparam>
<lparam>Address:820 2080</lparam>
<lparam>Address:821 2081</lparam>
<lparam>Address:822 2082</lparam>
<lparam>Address:823 2083</lparam>
<lparam>Address:824 2084</lparam>
<lparam>Address:825 2085</lparam>
<lparam>Address:826 2086</lparam>
<lparam>Address:827 2087</lparam>
<lparam>Address:828 2088</lparam>
<lparam>Address:829 2089</lparam>
<lparam>Address:830 2096</lparam>
<lparam>Address:831 2097</lparam>
<lparam>Address:832 2098</lparam>
<lparam>Address:833 2099</lparam>
<lparam>Address:834 2100</lparam>
<lparam>Address:835 2101</lparam>
<lparam>Address:836 2102</lparam>
<lparam>Address:837 2103</lparam>
<lparam>Address:838 2104</lparam>
<lparam>Address:839 2105</lparam>
<lparam>Address:840 2112</lparam>
<lparam>Address:841 2113</lparam>
<lparam>Address:842 2114</lparam>
<lparam>Address:843 2115</lparam>
<lparam>Address:844 2116</lparam>
<lparam>Address:845 2117</lparam>
<lparam>Address:846 2118</lparam>
<lparam>Address:847 2119</lparam>
<lparam>Address:848 2120</lparam>
<lparam>Address:849 2121</lparam>
<lparam>Address:850 2128</lparam>
<lparam>Address:851 2129</lparam>
<lparam>Address:852 2130</lparam>
<lparam>Address:853 2131</lparam>
<lparam>Address:854 2132</lparam>
<lparam>Address:855 2133</lparam>
<lparam>Address:856 2134</lparam>
<lparam>Address:857 2135</lparam>
<lparam>Address:858 2136</lparam>
<lparam>Address:859 2137</lparam>
<lparam>Address:860 2144</lparam>
<lparam>Address:861 2145</lparam>
<lparam>Address:862 2146</lparam>
<lparam>Address:863 2147</lparam>
<lparam>Address:864 2148</lparam>
<lparam>Address:865 2149</lparam>
<lparam>Address:866 2150</lparam>
<lparam>Address:867 2151</lparam>
<lparam>Address:868 2152</lparam>
<lparam>Address:869 2153</lparam>
<lparam>Address:870 2160</lparam>
<lparam>Address:871 2161</lparam>
<lparam>Address:872 2162</lparam>
<lparam>Address:873 2163</lparam>
<lparam>Address:874 2164</lparam>
<lparam>Address:875 2165</lparam>
<lparam>Address:876 2166</lparam>
<lparam>Address:877 2167</lparam>
<lparam>Address:878 2168</lparam>
<lparam>Address:879 2169</lparam>
<lparam>Address:880 2176</lparam>
<lparam>Address:881 2177</lparam>
<lparam>Address:882 2178</lparam>
<lparam>Address:883 2179</lparam>
<lparam>Address:884 2180</lparam>
<lparam>Address:885 2181</lparam>
<lparam>Address:886 2182</lparam>
<lparam>Address:887 2183</lparam>
<lparam>Address:888 2184</lparam>
<lparam>Address:889 2185</lparam>
<lparam>Address:890 2192</lparam>
<lparam>Address:891 2193</lparam>
<lparam>Address:892 2194</lparam>
<lparam>Address:893 2195</lparam>
<lparam>Address:894 2196</lparam>
<lparam>Address:895 2197</lparam>
<lparam>Address:896 2198</lparam>
<lparam>Address:897 2199</lparam>
<lparam>Address:898 2200</lparam>
<lparam>Address:899 2201</lparam>
<lparam>Address:900 2304</lparam>
<lparam>Address:901 2305</lparam>
<lparam>Address:902 2306</lparam>
<lparam>Address:903 2307</lparam>
<lparam>Address:904 2308</lparam>
<lparam>Address:905 2309</lparam>
<lparam>Address:906 2310</lparam>
<lparam>Address:907 2311</lparam>
<lparam>Address:908 2312</lparam>
<lparam>Address:909 2313</lparam>
<lparam>Address:910 2320</lparam>
<lparam>Address:911 2321</lparam>
<lparam>Address:912 2322</lparam>
<lparam>Address:913 2323</lparam>
<lparam>Address:914 2324</lparam>
<lparam>Address:915 2325</lparam>
<lparam>Address:916 2326</lparam>
<lparam>Address:917 2327</lparam>
<lparam>Address:918 2328</lparam>
<lparam>Address:919 2329</lparam>
<lparam>Address:920 2336</lparam>
<lparam>Address:921 2337</lparam>
<lparam>Address:922 2338</lparam>
<lparam>Address:923 2339</lparam>
<lparam>Address:924 2340</lparam>
<lparam>Address:925 2341</lparam>
<lparam>Address:926 2342</lparam>
<lparam>Address:927 2343</lparam>
<lparam>Address:928 2344</lparam>
<lparam>Address:929 2345</lparam>
<lparam>Address:930 2352</lparam>
<lparam>Address:931 2353</lparam>
<lparam>Address:932 2354</lparam>
<lparam>Address:933 2355</lparam>
<lparam>Address:934 2356</lparam>
<lparam>Address:935 2357</lparam>
<lparam>Address:936 2358</lparam>
<lparam>Address:937 2359</lparam>
<lparam>Address:938 2360</lparam>
<lparam>Address:939 2361</lparam>
<lparam>Address:940 2368</lparam>
<lparam>Address:941 2369</lparam>
<lparam>Address:942 2370</lparam>
<lparam>Address:943 2371</lparam>
<lparam>Address:944 2372</lparam>
<lparam>Address:945 2373</lparam>
<lparam>Address:946 2374</lparam>
<lparam>Address:947 2375</lparam>
<lparam>Address:948 2376</lparam>
<lparam>Address:949 2377</lparam>
<lparam>Address:950 2384</lparam>
<lparam>Address:951 2385</lparam>
<lparam>Address:952 2386</lparam>
<lparam>Address:953 2387</lparam>
<lparam>Address:954 2388</lparam>
<lparam>Address:955 2389</lparam>
<lparam>Address:956 2390</lparam>
<lparam>Address:957 2391</lparam>
<lparam>Address:958 2392</lparam>
<lparam>Address:959 2393</lparam>
<lparam>Address:960 2400</lparam>
<lparam>Address:961 2401</lparam>
<lparam>Address:962 2402</lparam>
<lparam>Address:963 2403</lparam>
<lparam>Address:964 2404</lparam>
<lparam>Address:965 2405</lparam>
<lparam>Address:966 2406</lparam>
<lparam>Address:967 2407</lparam>
<lparam>Address:968 2408</lparam>
<lparam>Address:969 2409</lparam>
<lparam>Address:970 2416</lparam>
<lparam>Address:971 2417</lparam>
<lparam>Address:972 2418</lparam>
<lparam>Address:973 2419</lparam>
<lparam>Address:974 2420</lparam>
<lparam>Address:975 2421</lparam>
<lparam>Address:976 2422</lparam>
<lparam>Address:977 2423</lparam>
<lparam>Address:978 2424</lparam>
<lparam>Address:979 2425</lparam>
<lparam>Address:980 2432</lparam>
<lparam>Address:981 2433</lparam>
<lparam>Address:982 2434</lparam>
<lparam>Address:983 2435</lparam>
<lparam>Address:984 2436</lparam>
<lparam>Address:985 2437</lparam>
<lparam>Address:986 2438</lparam>
<lparam>Address:987 2439</lparam>
<lparam>Address:988 2440</lparam>
<lparam>Address:989 2441</lparam>
<lparam>Address:990 2448</lparam>
<lparam>Address:991 2449</lparam>
<lparam>Address:992 2450</lparam>
<lparam>Address:993 2451</lparam>
<lparam>Address:994 2452</lparam>
<lparam>Address:995 2453</lparam>
<lparam>Address:996 2454</lparam>
<lparam>Address:997 2455</lparam>
<lparam>Address:998 2456</lparam>
<lparam>Address:999 2457</lparam>
<lparam>Address:1001 4097</lparam>
<lparam>Address:1002 4098</lparam>
<lparam>Address:1003 4099</lparam>
<lparam>Address:1004 4100</lparam>
<lparam>Address:1005 4101</lparam>
<lparam>Address:1006 4102</lparam>
<lparam>Address:1007 4103</lparam>
<lparam>Address:1008 4104</lparam>
<lparam>Address:1009 4105</lparam>
<lparam>Address:1010 4112</lparam>
<lparam>Address:1011 4113</lparam>
<lparam>Address:1012 4114</lparam>
<lparam>Address:1013 4115</lparam>
<lparam>Address:1014 4116</lparam>
<lparam>Address:1015 4117</lparam>
<lparam>Address:1016 4118</lparam>
<lparam>Address:1017 4119</lparam>
<lparam>Address:1018 4120</lparam>
<lparam>Address:1019 4121</lparam>
<lparam>Address:1020 4128</lparam>
<lparam>Address:1021 4129</lparam>
<lparam>Address:1022 4130</lparam>
<lparam>Address:1023 4131</lparam>
<lparam>Address:1024 4132</lparam>
<lparam>Address:1025 4133</lparam>
<lparam>Address:1026 4134</lparam>
<lparam>Address:1027 4135</lparam>
<lparam>Address:1028 4136</lparam>
<lparam>Address:1029 4137</lparam>
<lparam>Address:1030 4144</lparam>
<lparam>Address:1031 4145</lparam>
<lparam>Address:1032 4146</lparam>
<lparam>Address:1033 4147</lparam>
<lparam>Address:1034 4148</lparam>
<lparam>Address:1035 4149</lparam>
<lparam>Address:1036 4150</lparam>
<lparam>Address:1037 4151</lparam>
<lparam>Address:1038 4152</lparam>
<lparam>Address:1039 4153</lparam>
<lparam>Address:1040 4160</lparam>
<lparam>Address:1041 4161</lparam>
<lparam>Address:1042 4162</lparam>
<lparam>Address:1043 4163</lparam>
<lparam>Address:1044 4164</lparam>
<lparam>Address:1045 4165</lparam>
<lparam>Address:1046 4166</lparam>
<lparam>Address:1047 4167</lparam>
<lparam>Address:1048 4168</lparam>
<lparam>Address:1049 4169</lparam>
<lparam>Address:1050 4176</lparam>
<lparam>Address:1051 4177</lparam>
<lparam>Address:1052 4178</lparam>
<lparam>Address:1053 4179</lparam>
<lparam>Address:1054 4180</lparam>
<lparam>Address:1055 4181</lparam>
<lparam>Address:1056 4182</lparam>
<lparam>Address:1057 4183</lparam>
<lparam>Address:1058 4184</lparam>
<lparam>Address:1059 4185</lparam>
<lparam>Address:1060 4192</lparam>
<lparam>Address:1061 4193</lparam>
<lparam>Address:1062 4194</lparam>
<lparam>Address:1063 4195</lparam>
<lparam>Address:1064 4196</lparam>
<lparam>Address:1065 4197</lparam>
<lparam>Address:1066 4198</lparam>
<lparam>Address:1067 4199</lparam>
<lparam>Address:1068 4200</lparam>
<lparam>Address:1069 4201</lparam>
<lparam>Address:1070 4208</lparam>
<lparam>Address:1071 4209</lparam>
<lparam>Address:1072 4210</lparam>
<lparam>Address:1073 4211</lparam>
<lparam>Address:1074 4212</lparam>
<lparam>Address:1075 4213</lparam>
<lparam>Address:1076 4214</lparam>
<lparam>Address:1077 4215</lparam>
<lparam>Address:1078 4216</lparam>
<lparam>Address:1079 4217</lparam>
<lparam>Address:1080 4224</lparam>
<lparam>Address:1081 4225</lparam>
<lparam>Address:1082 4226</lparam>
<lparam>Address:1083 4227</lparam>
<lparam>Address:1084 4228</lparam>
<lparam>Address:1085 4229</lparam>
<lparam>Address:1086 4230</lparam>
<lparam>Address:1087 4231</lparam>
<lparam>Address:1088 4232</lparam>
<lparam>Address:1089 4233</lparam>
<lparam>Address:1090 4240</lparam>
<lparam>Address:1091 4241</lparam>
<lparam>Address:1092 4242</lparam>
<lparam>Address:1093 4243</lparam>
<lparam>Address:1094 4244</lparam>
<lparam>Address:1095 4245</lparam>
<lparam>Address:1096 4246</lparam>
<lparam>Address:1097 4247</lparam>
<lparam>Address:1098 4248</lparam>
<lparam>Address:1099 4249</lparam>
<lparam>Address:1100 4352</lparam>
<lparam>Address:1101 4353</lparam>
<lparam>Address:1102 4354</lparam>
<lparam>Address:1103 4355</lparam>
<lparam>Address:1104 4356</lparam>
<lparam>Address:1105 4357</lparam>
<lparam>Address:1106 4358</lparam>
<lparam>Address:1107 4359</lparam>
<lparam>Address:1108 4360</lparam>
<lparam>Address:1109 4361</lparam>
<lparam>Address:1110 4368</lparam>
<lparam>Address:1111 4369</lparam>
<lparam>Address:1112 4370</lparam>
<lparam>Address:1113 4371</lparam>
<lparam>Address:1114 4372</lparam>
<lparam>Address:1115 4373</lparam>
<lparam>Address:1116 4374</lparam>
<lparam>Address:1117 4375</lparam>
<lparam>Address:1118 4376</lparam>
<lparam>Address:1119 4377</lparam>
<lparam>Address:1120 4384</lparam>
<lparam>Address:1121 4385</lparam>
<lparam>Address:1122 4386</lparam>
<lparam>Address:1123 4387</lparam>
<lparam>Address:1124 4388</lparam>
<lparam>Address:1125 4389</lparam>
<lparam>Address:1126 4390</lparam>
<lparam>Address:1127 4391</lparam>
<lparam>Address:1128 4392</lparam>
<lparam>Address:1129 4393</lparam>
<lparam>Address:1130 4400</lparam>
<lparam>Address:1131 4401</lparam>
<lparam>Address:1132 4402</lparam>
<lparam>Address:1133 4403</lparam>
<lparam>Address:1134 4404</lparam>
<lparam>Address:1135 4405</lparam>
<lparam>Address:1136 4406</lparam>
<lparam>Address:1137 4407</lparam>
<lparam>Address:1138 4408</lparam>
<lparam>Address:1139 4409</lparam>
<lparam>Address:1140 4416</lparam>
<lparam>Address:1141 4417</lparam>
<lparam>Address:1142 4418</lparam>
<lparam>Address:1143 4419</lparam>
<lparam>Address:1144 4420</lparam>
<lparam>Address:1145 4421</lparam>
<lparam>Address:1146 4422</lparam>
<lparam>Address:1147 4423</lparam>
<lparam>Address:1148 4424</lparam>
<lparam>Address:1149 4425</lparam>
<lparam>Address:1150 4432</lparam>
<lparam>Address:1151 4433</lparam>
<lparam>Address:1152 4434</lparam>
<lparam>Address:1153 4435</lparam>
<lparam>Address:1154 4436</lparam>
<lparam>Address:1155 4437</lparam>
<lparam>Address:1156 4438</lparam>
<lparam>Address:1157 4439</lparam>
<lparam>Address:1158 4440</lparam>
<lparam>Address:1159 4441</lparam>
<lparam>Address:1160 4448</lparam>
<lparam>Address:1161 4449</lparam>
<lparam>Address:1162 4450</lparam>
<lparam>Address:1163 4451</lparam>
<lparam>Address:1164 4452</lparam>
<lparam>Address:1165 4453</lparam>
<lparam>Address:1166 4454</lparam>
<lparam>Address:1167 4455</lparam>
<lparam>Address:1168 4456</lparam>
<lparam>Address:1169 4457</lparam>
<lparam>Address:1170 4464</lparam>
<lparam>Address:1171 4465</lparam>
<lparam>Address:1172 4466</lparam>
<lparam>Address:1173 4467</lparam>
<lparam>Address:1174 4468</lparam>
<lparam>Address:1175 4469</lparam>
<lparam>Address:1176 4470</lparam>
<lparam>Address:1177 4471</lparam>
<lparam>Address:1178 4472</lparam>
<lparam>Address:1179 4473</lparam>
<lparam>Address:1180 4480</lparam>
<lparam>Address:1181 4481</lparam>
<lparam>Address:1182 4482</lparam>
<lparam>Address:1183 4483</lparam>
<lparam>Address:1184 4484</lparam>
<lparam>Address:1185 4485</lparam>
<lparam>Address:1186 4486</lparam>
<lparam>Address:1187 4487</lparam>
<lparam>Address:1188 4488</lparam>
<lparam>Address:1189 4489</lparam>
<lparam>Address:1190 4496</lparam>
<lparam>Address:1191 4497</lparam>
<lparam>Address:1192 4498</lparam>
<lparam>Address:1193 4499</lparam>
<lparam>Address:1194 4500</lparam>
<lparam>Address:1195 4501</lparam>
<lparam>Address:1196 4502</lparam>
<lparam>Address:1197 4503</lparam>
<lparam>Address:1198 4504</lparam>
<lparam>Address:1199 4505</lparam>
<lparam>Address:1200 4608</lparam>
<lparam>Address:1201 4609</lparam>
<lparam>Address:1202 4610</lparam>
<lparam>Address:1203 4611</lparam>
<lparam>Address:1204 4612</lparam>
<lparam>Address:1205 4613</lparam>
<lparam>Address:1206 4614</lparam>
<lparam>Address:1207 4615</lparam>
<lparam>Address:1208 4616</lparam>
<lparam>Address:1209 4617</lparam>
<lparam>Address:1210 4624</lparam>
<lparam>Address:1211 4625</lparam>
<lparam>Address:1212 4626</lparam>
<lparam>Address:1213 4627</lparam>
<lparam>Address:1214 4628</lparam>
<lparam>Address:1215 4629</lparam>
<lparam>Address:1216 4630</lparam>
<lparam>Address:1217 4631</lparam>
<lparam>Address:1218 4632</lparam>
<lparam>Address:1219 4633</lparam>
<lparam>Address:1220 4640</lparam>
<lparam>Address:1221 4641</lparam>
<lparam>Address:1222 4642</lparam>
<lparam>Address:1223 4643</lparam>
<lparam>Address:1224 4644</lparam>
<lparam>Address:1225 4645</lparam>
<lparam>Address:1226 4646</lparam>
<lparam>Address:1227 4647</lparam>
<lparam>Address:1228 4648</lparam>
<lparam>Address:1229 4649</lparam>
<lparam>Address:1230 4656</lparam>
<lparam>Address:1231 4657</lparam>
<lparam>Address:1232 4658</lparam>
<lparam>Address:1233 4659</lparam>
<lparam>Address:1234 4660</lparam>
<lparam>Address:1235 4661</lparam>
<lparam>Address:1236 4662</lparam>
<lparam>Address:1237 4663</lparam>
<lparam>Address:1238 4664</lparam>
<lparam>Address:1239 4665</lparam>
<lparam>Address:1240 4672</lparam>
<lparam>Address:1241 4673</lparam>
<lparam>Address:1242 4674</lparam>
<lparam>Address:1243 4675</lparam>
<lparam>Address:1244 4676</lparam>
<lparam>Address:1245 4677</lparam>
<lparam>Address:1246 4678</lparam>
<lparam>Address:1247 4679</lparam>
<lparam>Address:1248 4680</lparam>
<lparam>Address:1249 4681</lparam>
<lparam>Address:1250 4688</lparam>
<lparam>Address:1251 4689</lparam>
<lparam>Address:1252 4690</lparam>
<lparam>Address:1253 4691</lparam>
<lparam>Address:1254 4692</lparam>
<lparam>Address:1255 4693</lparam>
<lparam>Address:1256 4694</lparam>
<lparam>Address:1257 4695</lparam>
<lparam>Address:1258 4696</lparam>
<lparam>Address:1259 4697</lparam>
<lparam>Address:1260 4704</lparam>
<lparam>Address:1261 4705</lparam>
<lparam>Address:1262 4706</lparam>
<lparam>Address:1263 4707</lparam>
<lparam>Address:1264 4708</lparam>
<lparam>Address:1265 4709</lparam>
<lparam>Address:1266 4710</lparam>
<lparam>Address:1267 4711</lparam>
<lparam>Address:1268 4712</lparam>
<lparam>Address:1269 4713</lparam>
<lparam>Address:1270 4720</lparam>
<lparam>Address:1271 4721</lparam>
<lparam>Address:1272 4722</lparam>
<lparam>Address:1273 4723</lparam>
<lparam>Address:1274 4724</lparam>
<lparam>Address:1275 4725</lparam>
<lparam>Address:1276 4726</lparam>
<lparam>Address:1277 4727</lparam>
<lparam>Address:1278 4728</lparam>
<lparam>Address:1279 4729</lparam>
<lparam>Address:1280 4736</lparam>
<lparam>Address:1281 4737</lparam>
<lparam>Address:1282 4738</lparam>
<lparam>Address:1283 4739</lparam>
<lparam>Address:1284 4740</lparam>
<lparam>Address:1285 4741</lparam>
<lparam>Address:1286 4742</lparam>
<lparam>Address:1287 4743</lparam>
<lparam>Address:1288 4744</lparam>
<lparam>Address:1289 4745</lparam>
<lparam>Address:1290 4752</lparam>
<lparam>Address:1291 4753</lparam>
<lparam>Address:1292 4754</lparam>
<lparam>Address:1293 4755</lparam>
<lparam>Address:1294 4756</lparam>
<lparam>Address:1295 4757</lparam>
<lparam>Address:1296 4758</lparam>
<lparam>Address:1297 4759</lparam>
<lparam>Address:1298 4760</lparam>
<lparam>Address:1299 4761</lparam>
<lparam>Address:1300 4864</lparam>
<lparam>Address:1301 4865</lparam>
<lparam>Address:1302 4866</lparam>
<lparam>Address:1303 4867</lparam>
<lparam>Address:1304 4868</lparam>
<lparam>Address:1305 4869</lparam>
<lparam>Address:1306 4870</lparam>
<lparam>Address:1307 4871</lparam>
<lparam>Address:1308 4872</lparam>
<lparam>Address:1309 4873</lparam>
<lparam>Address:1310 4880</lparam>
<lparam>Address:1311 4881</lparam>
<lparam>Address:1312 4882</lparam>
<lparam>Address:1313 4883</lparam>
<lparam>Address:1314 4884</lparam>
<lparam>Address:1315 4885</lparam>
<lparam>Address:1316 4886</lparam>
<lparam>Address:1317 4887</lparam>
<lparam>Address:1318 4888</lparam>
<lparam>Address:1319 4889</lparam>
<lparam>Address:1320 4896</lparam>
<lparam>Address:1321 4897</lparam>
<lparam>Address:1322 4898</lparam>
<lparam>Address:1323 4899</lparam>
<lparam>Address:1324 4900</lparam>
<lparam>Address:1325 4901</lparam>
<lparam>Address:1326 4902</lparam>
<lparam>Address:1327 4903</lparam>
<lparam>Address:1328 4904</lparam>
<lparam>Address:1329 4905</lparam>
<lparam>Address:1330 4912</lparam>
<lparam>Address:1331 4913</lparam>
<lparam>Address:1332 4914</lparam>
<lparam>Address:1333 4915</lparam>
<lparam>Address:1334 4916</lparam>
<lparam>Address:1335 4917</lparam>
<lparam>Address:1336 4918</lparam>
<lparam>Address:1337 4919</lparam>
<lparam>Address:1338 4920</lparam>
<lparam>Address:1339 4921</lparam>
<lparam>Address:1340 4928</lparam>
<lparam>Address:1341 4929</lparam>
<lparam>Address:1342 4930</lparam>
<lparam>Address:1343 4931</lparam>
<lparam>Address:1344 4932</lparam>
<lparam>Address:1345 4933</lparam>
<lparam>Address:1346 4934</lparam>
<lparam>Address:1347 4935</lparam>
<lparam>Address:1348 4936</lparam>
<lparam>Address:1349 4937</lparam>
<lparam>Address:1350 4944</lparam>
<lparam>Address:1351 4945</lparam>
<lparam>Address:1352 4946</lparam>
<lparam>Address:1353 4947</lparam>
<lparam>Address:1354 4948</lparam>
<lparam>Address:1355 4949</lparam>
<lparam>Address:1356 4950</lparam>
<lparam>Address:1357 4951</lparam>
<lparam>Address:1358 4952</lparam>
<lparam>Address:1359 4953</lparam>
<lparam>Address:1360 4960</lparam>
<lparam>Address:1361 4961</lparam>
<lparam>Address:1362 4962</lparam>
<lparam>Address:1363 4963</lparam>
<lparam>Address:1364 4964</lparam>
<lparam>Address:1365 4965</lparam>
<lparam>Address:1366 4966</lparam>
<lparam>Address:1367 4967</lparam>
<lparam>Address:1368 4968</lparam>
<lparam>Address:1369 4969</lparam>
<lparam>Address:1370 4976</lparam>
<lparam>Address:1371 4977</lparam>
<lparam>Address:1372 4978</lparam>
<lparam>Address:1373 4979</lparam>
<lparam>Address:1374 4980</lparam>
<lparam>Address:1375 4981</lparam>
<lparam>Address:1376 4982</lparam>
<lparam>Address:1377 4983</lparam>
<lparam>Address:1378 4984</lparam>
<lparam>Address:1379 4985</lparam>
<lparam>Address:1380 4992</lparam>
<lparam>Address:1381 4993</lparam>
<lparam>Address:1382 4994</lparam>
<lparam>Address:1383 4995</lparam>
<lparam>Address:1384 4996</lparam>
<lparam>Address:1385 4997</lparam>
<lparam>Address:1386 4998</lparam>
<lparam>Address:1387 4999</lparam>
<lparam>Address:1388 5000</lparam>
<lparam>Address:1389 5001</lparam>
<lparam>Address:1390 5008</lparam>
<lparam>Address:1391 5009</lparam>
<lparam>Address:1392 5010</lparam>
<lparam>Address:1393 5011</lparam>
<lparam>Address:1394 5012</lparam>
<lparam>Address:1395 5013</lparam>
<lparam>Address:1396 5014</lparam>
<lparam>Address:1397 5015</lparam>
<lparam>Address:1398 5016</lparam>
<lparam>Address:1399 5017</lparam>
<lparam>Address:1400 5120</lparam>
<lparam>Address:1401 5121</lparam>
<lparam>Address:1402 5122</lparam>
<lparam>Address:1403 5123</lparam>
<lparam>Address:1404 5124</lparam>
<lparam>Address:1405 5125</lparam>
<lparam>Address:1406 5126</lparam>
<lparam>Address:1407 5127</lparam>
<lparam>Address:1408 5128</lparam>
<lparam>Address:1409 5129</lparam>
<lparam>Address:1410 5136</lparam>
<lparam>Address:1411 5137</lparam>
<lparam>Address:1412 5138</lparam>
<lparam>Address:1413 5139</lparam>
<lparam>Address:1414 5140</lparam>
<lparam>Address:1415 5141</lparam>
<lparam>Address:1416 5142</lparam>
<lparam>Address:1417 5143</lparam>
<lparam>Address:1418 5144</lparam>
<lparam>Address:1419 5145</lparam>
<lparam>Address:1420 5152</lparam>
<lparam>Address:1421 5153</lparam>
<lparam>Address:1422 5154</lparam>
<lparam>Address:1423 5155</lparam>
<lparam>Address:1424 5156</lparam>
<lparam>Address:1425 5157</lparam>
<lparam>Address:1426 5158</lparam>
<lparam>Address:1427 5159</lparam>
<lparam>Address:1428 5160</lparam>
<lparam>Address:1429 5161</lparam>
<lparam>Address:1430 5168</lparam>
<lparam>Address:1431 5169</lparam>
<lparam>Address:1432 5170</lparam>
<lparam>Address:1433 5171</lparam>
<lparam>Address:1434 5172</lparam>
<lparam>Address:1435 5173</lparam>
<lparam>Address:1436 5174</lparam>
<lparam>Address:1437 5175</lparam>
<lparam>Address:1438 5176</lparam>
<lparam>Address:1439 5177</lparam>
<lparam>Address:1440 5184</lparam>
<lparam>Address:1441 5185</lparam>
<lparam>Address:1442 5186</lparam>
<lparam>Address:1443 5187</lparam>
<lparam>Address:1444 5188</lparam>
<lparam>Address:1445 5189</lparam>
<lparam>Address:1446 5190</lparam>
<lparam>Address:1447 5191</lparam>
<lparam>Address:1448 5192</lparam>
<lparam>Address:1449 5193</lparam>
<lparam>Address:1450 5200</lparam>
<lparam>Address:1451 5201</lparam>
<lparam>Address:1452 5202</lparam>
<lparam>Address:1453 5203</lparam>
<lparam>Address:1454 5204</lparam>
<lparam>Address:1455 5205</lparam>
<lparam>Address:1456 5206</lparam>
<lparam>Address:1457 5207</lparam>
<lparam>Address:1458 5208</lparam>
<lparam>Address:1459 5209</lparam>
<lparam>Address:1460 5216</lparam>
<lparam>Address:1461 5217</lparam>
<lparam>Address:1462 5218</lparam>
<lparam>Address:1463 5219</lparam>
<lparam>Address:1464 5220</lparam>
<lparam>Address:1465 5221</lparam>
<lparam>Address:1466 5222</lparam>
<lparam>Address:1467 5223</lparam>
<lparam>Address:1468 5224</lparam>
<lparam>Address:1469 5225</lparam>
<lparam>Address:1470 5232</lparam>
<lparam>Address:1471 5233</lparam>
<lparam>Address:1472 5234</lparam>
<lparam>Address:1473 5235</lparam>
<lparam>Address:1474 5236</lparam>
<lparam>Address:1475 5237</lparam>
<lparam>Address:1476 5238</lparam>
<lparam>Address:1477 5239</lparam>
<lparam>Address:1478 5240</lparam>
<lparam>Address:1479 5241</lparam>
<lparam>Address:1480 5248</lparam>
<lparam>Address:1481 5249</lparam>
<lparam>Address:1482 5250</lparam>
<lparam>Address:1483 5251</lparam>
<lparam>Address:1484 5252</lparam>
<lparam>Address:1485 5253</lparam>
<lparam>Address:1486 5254</lparam>
<lparam>Address:1487 5255</lparam>
<lparam>Address:1488 5256</lparam>
<lparam>Address:1489 5257</lparam>
<lparam>Address:1490 5264</lparam>
<lparam>Address:1491 5265</lparam>
<lparam>Address:1492 5266</lparam>
<lparam>Address:1493 5267</lparam>
<lparam>Address:1494 5268</lparam>
<lparam>Address:1495 5269</lparam>
<lparam>Address:1496 5270</lparam>
<lparam>Address:1497 5271</lparam>
<lparam>Address:1498 5272</lparam>
<lparam>Address:1499 5273</lparam>
<lparam>Address:1500 5376</lparam>
<lparam>Address:1501 5377</lparam>
<lparam>Address:1502 5378</lparam>
<lparam>Address:1503 5379</lparam>
<lparam>Address:1504 5380</lparam>
<lparam>Address:1505 5381</lparam>
<lparam>Address:1506 5382</lparam>
<lparam>Address:1507 5383</lparam>
<lparam>Address:1508 5384</lparam>
<lparam>Address:1509 5385</lparam>
<lparam>Address:1510 5392</lparam>
<lparam>Address:1511 5393</lparam>
<lparam>Address:1512 5394</lparam>
<lparam>Address:1513 5395</lparam>
<lparam>Address:1514 5396</lparam>
<lparam>Address:1515 5397</lparam>
<lparam>Address:1516 5398</lparam>
<lparam>Address:1517 5399</lparam>
<lparam>Address:1518 5400</lparam>
<lparam>Address:1519 5401</lparam>
<lparam>Address:1520 5408</lparam>
<lparam>Address:1521 5409</lparam>
<lparam>Address:1522 5410</lparam>
<lparam>Address:1523 5411</lparam>
<lparam>Address:1524 5412</lparam>
<lparam>Address:1525 5413</lparam>
<lparam>Address:1526 5414</lparam>
<lparam>Address:1527 5415</lparam>
<lparam>Address:1528 5416</lparam>
<lparam>Address:1529 5417</lparam>
<lparam>Address:1530 5424</lparam>
<lparam>Address:1531 5425</lparam>
<lparam>Address:1532 5426</lparam>
<lparam>Address:1533 5427</lparam>
<lparam>Address:1534 5428</lparam>
<lparam>Address:1535 5429</lparam>
<lparam>Address:1536 5430</lparam>
<lparam>Address:1537 5431</lparam>
<lparam>Address:1538 5432</lparam>
<lparam>Address:1539 5433</lparam>
<lparam>Address:1540 5440</lparam>
<lparam>Address:1541 5441</lparam>
<lparam>Address:1542 5442</lparam>
<lparam>Address:1543 5443</lparam>
<lparam>Address:1544 5444</lparam>
<lparam>Address:1545 5445</lparam>
<lparam>Address:1546 5446</lparam>
<lparam>Address:1547 5447</lparam>
<lparam>Address:1548 5448</lparam>
<lparam>Address:1549 5449</lparam>
<lparam>Address:1550 5456</lparam>
<lparam>Address:1551 5457</lparam>
<lparam>Address:1552 5458</lparam>
<lparam>Address:1553 5459</lparam>
<lparam>Address:1554 5460</lparam>
<lparam>Address:1555 5461</lparam>
<lparam>Address:1556 5462</lparam>
<lparam>Address:1557 5463</lparam>
<lparam>Address:1558 5464</lparam>
<lparam>Address:1559 5465</lparam>
<lparam>Address:1560 5472</lparam>
<lparam>Address:1561 5473</lparam>
<lparam>Address:1562 5474</lparam>
<lparam>Address:1563 5475</lparam>
<lparam>Address:1564 5476</lparam>
<lparam>Address:1565 5477</lparam>
<lparam>Address:1566 5478</lparam>
<lparam>Address:1567 5479</lparam>
<lparam>Address:1568 5480</lparam>
<lparam>Address:1569 5481</lparam>
<lparam>Address:1570 5488</lparam>
<lparam>Address:1571 5489</lparam>
<lparam>Address:1572 5490</lparam>
<lparam>Address:1573 5491</lparam>
<lparam>Address:1574 5492</lparam>
<lparam>Address:1575 5493</lparam>
<lparam>Address:1576 5494</lparam>
<lparam>Address:1577 5495</lparam>
<lparam>Address:1578 5496</lparam>
<lparam>Address:1579 5497</lparam>
<lparam>Address:1580 5504</lparam>
<lparam>Address:1581 5505</lparam>
<lparam>Address:1582 5506</lparam>
<lparam>Address:1583 5507</lparam>
<lparam>Address:1584 5508</lparam>
<lparam>Address:1585 5509</lparam>
<lparam>Address:1586 5510</lparam>
<lparam>Address:1587 5511</lparam>
<lparam>Address:1588 5512</lparam>
<lparam>Address:1589 5513</lparam>
<lparam>Address:1590 5520</lparam>
<lparam>Address:1591 5521</lparam>
<lparam>Address:1592 5522</lparam>
<lparam>Address:1593 5523</lparam>
<lparam>Address:1594 5524</lparam>
<lparam>Address:1595 5525</lparam>
<lparam>Address:1596 5526</lparam>
<lparam>Address:1597 5527</lparam>
<lparam>Address:1598 5528</lparam>
<lparam>Address:1599 5529</lparam>
<lparam>Address:1600 5632</lparam>
<lparam>Address:1601 5633</lparam>
<lparam>Address:1602 5634</lparam>
<lparam>Address:1603 5635</lparam>
<lparam>Address:1604 5636</lparam>
<lparam>Address:1605 5637</lparam>
<lparam>Address:1606 5638</lparam>
<lparam>Address:1607 5639</lparam>
<lparam>Address:1608 5640</lparam>
<lparam>Address:1609 5641</lparam>
<lparam>Address:1610 5648</lparam>
<lparam>Address:1611 5649</lparam>
<lparam>Address:1612 5650</lparam>
<lparam>Address:1613 5651</lparam>
<lparam>Address:1614 5652</lparam>
<lparam>Address:1615 5653</lparam>
<lparam>Address:1616 5654</lparam>
<lparam>Address:1617 5655</lparam>
<lparam>Address:1618 5656</lparam>
<lparam>Address:1619 5657</lparam>
<lparam>Address:1620 5664</lparam>
<lparam>Address:1621 5665</lparam>
<lparam>Address:1622 5666</lparam>
<lparam>Address:1623 5667</lparam>
<lparam>Address:1624 5668</lparam>
<lparam>Address:1625 5669</lparam>
<lparam>Address:1626 5670</lparam>
<lparam>Address:1627 5671</lparam>
<lparam>Address:1628 5672</lparam>
<lparam>Address:1629 5673</lparam>
<lparam>Address:1630 5680</lparam>
<lparam>Address:1631 5681</lparam>
<lparam>Address:1632 5682</lparam>
<lparam>Address:1633 5683</lparam>
<lparam>Address:1634 5684</lparam>
<lparam>Address:1635 5685</lparam>
<lparam>Address:1636 5686</lparam>
<lparam>Address:1637 5687</lparam>
<lparam>Address:1638 5688</lparam>
<lparam>Address:1639 5689</lparam>
<lparam>Address:1640 5696</lparam>
<lparam>Address:1641 5697</lparam>
<lparam>Address:1642 5698</lparam>
<lparam>Address:1643 5699</lparam>
<lparam>Address:1644 5700</lparam>
<lparam>Address:1645 5701</lparam>
<lparam>Address:1646 5702</lparam>
<lparam>Address:1647 5703</lparam>
<lparam>Address:1648 5704</lparam>
<lparam>Address:1649 5705</lparam>
<lparam>Address:1650 5712</lparam>
<lparam>Address:1651 5713</lparam>
<lparam>Address:1652 5714</lparam>
<lparam>Address:1653 5715</lparam>
<lparam>Address:1654 5716</lparam>
<lparam>Address:1655 5717</lparam>
<lparam>Address:1656 5718</lparam>
<lparam>Address:1657 5719</lparam>
<lparam>Address:1658 5720</lparam>
<lparam>Address:1659 5721</lparam>
<lparam>Address:1660 5728</lparam>
<lparam>Address:1661 5729</lparam>
<lparam>Address:1662 5730</lparam>
<lparam>Address:1663 5731</lparam>
<lparam>Address:1664 5732</lparam>
<lparam>Address:1665 5733</lparam>
<lparam>Address:1666 5734</lparam>
<lparam>Address:1667 5735</lparam>
<lparam>Address:1668 5736</lparam>
<lparam>Address:1669 5737</lparam>
<lparam>Address:1670 5744</lparam>
<lparam>Address:1671 5745</lparam>
<lparam>Address:1672 5746</lparam>
<lparam>Address:1673 5747</lparam>
<lparam>Address:1674 5748</lparam>
<lparam>Address:1675 5749</lparam>
<lparam>Address:1676 5750</lparam>
<lparam>Address:1677 5751</lparam>
<lparam>Address:1678 5752</lparam>
<lparam>Address:1679 5753</lparam>
<lparam>Address:1680 5760</lparam>
<lparam>Address:1681 5761</lparam>
<lparam>Address:1682 5762</lparam>
<lparam>Address:1683 5763</lparam>
<lparam>Address:1684 5764</lparam>
<lparam>Address:1685 5765</lparam>
<lparam>Address:1686 5766</lparam>
<lparam>Address:1687 5767</lparam>
<lparam>Address:1688 5768</lparam>
<lparam>Address:1689 5769</lparam>
<lparam>Address:1690 5776</lparam>
<lparam>Address:1691 5777</lparam>
<lparam>Address:1692 5778</lparam>
<lparam>Address:1693 5779</lparam>
<lparam>Address:1694 5780</lparam>
<lparam>Address:1695 5781</lparam>
<lparam>Address:1696 5782</lparam>
<lparam>Address:1697 5783</lparam>
<lparam>Address:1698 5784</lparam>
<lparam>Address:1699 5785</lparam>
<lparam>Address:1700 5888</lparam>
<lparam>Address:1701 5889</lparam>
<lparam>Address:1702 5890</lparam>
<lparam>Address:1703 5891</lparam>
<lparam>Address:1704 5892</lparam>
<lparam>Address:1705 5893</lparam>
<lparam>Address:1706 5894</lparam>
<lparam>Address:1707 5895</lparam>
<lparam>Address:1708 5896</lparam>
<lparam>Address:1709 5897</lparam>
<lparam>Address:1710 5904</lparam>
<lparam>Address:1711 5905</lparam>
<lparam>Address:1712 5906</lparam>
<lparam>Address:1713 5907</lparam>
<lparam>Address:1714 5908</lparam>
<lparam>Address:1715 5909</lparam>
<lparam>Address:1716 5910</lparam>
<lparam>Address:1717 5911</lparam>
<lparam>Address:1718 5912</lparam>
<lparam>Address:1719 5913</lparam>
<lparam>Address:1720 5920</lparam>
<lparam>Address:1721 5921</lparam>
<lparam>Address:1722 5922</lparam>
<lparam>Address:1723 5923</lparam>
<lparam>Address:1724 5924</lparam>
<lparam>Address:1725 5925</lparam>
<lparam>Address:1726 5926</lparam>
<lparam>Address:1727 5927</lparam>
<lparam>Address:1728 5928</lparam>
<lparam>Address:1729 5929</lparam>
<lparam>Address:1730 5936</lparam>
<lparam>Address:1731 5937</lparam>
<lparam>Address:1732 5938</lparam>
<lparam>Address:1733 5939</lparam>
<lparam>Address:1734 5940</lparam>
<lparam>Address:1735 5941</lparam>
<lparam>Address:1736 5942</lparam>
<lparam>Address:1737 5943</lparam>
<lparam>Address:1738 5944</lparam>
<lparam>Address:1739 5945</lparam>
<lparam>Address:1740 5952</lparam>
<lparam>Address:1741 5953</lparam>
<lparam>Address:1742 5954</lparam>
<lparam>Address:1743 5955</lparam>
<lparam>Address:1744 5956</lparam>
<lparam>Address:1745 5957</lparam>
<lparam>Address:1746 5958</lparam>
<lparam>Address:1747 5959</lparam>
<lparam>Address:1748 5960</lparam>
<lparam>Address:1749 5961</lparam>
<lparam>Address:1750 5968</lparam>
<lparam>Address:1751 5969</lparam>
<lparam>Address:1752 5970</lparam>
<lparam>Address:1753 5971</lparam>
<lparam>Address:1754 5972</lparam>
<lparam>Address:1755 5973</lparam>
<lparam>Address:1756 5974</lparam>
<lparam>Address:1757 5975</lparam>
<lparam>Address:1758 5976</lparam>
<lparam>Address:1759 5977</lparam>
<lparam>Address:1760 5984</lparam>
<lparam>Address:1761 5985</lparam>
<lparam>Address:1762 5986</lparam>
<lparam>Address:1763 5987</lparam>
<lparam>Address:1764 5988</lparam>
<lparam>Address:1765 5989</lparam>
<lparam>Address:1766 5990</lparam>
<lparam>Address:1767 5991</lparam>
<lparam>Address:1768 5992</lparam>
<lparam>Address:1769 5993</lparam>
<lparam>Address:1770 6000</lparam>
<lparam>Address:1771 6001</lparam>
<lparam>Address:1772 6002</lparam>
<lparam>Address:1773 6003</lparam>
<lparam>Address:1774 6004</lparam>
<lparam>Address:1775 6005</lparam>
<lparam>Address:1776 6006</lparam>
<lparam>Address:1777 6007</lparam>
<lparam>Address:1778 6008</lparam>
<lparam>Address:1779 6009</lparam>
<lparam>Address:1780 6016</lparam>
<lparam>Address:1781 6017</lparam>
<lparam>Address:1782 6018</lparam>
<lparam>Address:1783 6019</lparam>
<lparam>Address:1784 6020</lparam>
<lparam>Address:1785 6021</lparam>
<lparam>Address:1786 6022</lparam>
<lparam>Address:1787 6023</lparam>
<lparam>Address:1788 6024</lparam>
<lparam>Address:1789 6025</lparam>
<lparam>Address:1790 6032</lparam>
<lparam>Address:1791 6033</lparam>
<lparam>Address:1792 6034</lparam>
<lparam>Address:1793 6035</lparam>
<lparam>Address:1794 6036</lparam>
<lparam>Address:1795 6037</lparam>
<lparam>Address:1796 6038</lparam>
<lparam>Address:1797 6039</lparam>
<lparam>Address:1798 6040</lparam>
<lparam>Address:1799 6041</lparam>
<lparam>Address:1800 6144</lparam>
<lparam>Address:1801 6145</lparam>
<lparam>Address:1802 6146</lparam>
<lparam>Address:1803 6147</lparam>
<lparam>Address:1804 6148</lparam>
<lparam>Address:1805 6149</lparam>
<lparam>Address:1806 6150</lparam>
<lparam>Address:1807 6151</lparam>
<lparam>Address:1808 6152</lparam>
<lparam>Address:1809 6153</lparam>
<lparam>Address:1810 6160</lparam>
<lparam>Address:1811 6161</lparam>
<lparam>Address:1812 6162</lparam>
<lparam>Address:1813 6163</lparam>
<lparam>Address:1814 6164</lparam>
<lparam>Address:1815 6165</lparam>
<lparam>Address:1816 6166</lparam>
<lparam>Address:1817 6167</lparam>
<lparam>Address:1818 6168</lparam>
<lparam>Address:1819 6169</lparam>
<lparam>Address:1820 6176</lparam>
<lparam>Address:1821 6177</lparam>
<lparam>Address:1822 6178</lparam>
<lparam>Address:1823 6179</lparam>
<lparam>Address:1824 6180</lparam>
<lparam>Address:1825 6181</lparam>
<lparam>Address:1826 6182</lparam>
<lparam>Address:1827 6183</lparam>
<lparam>Address:1828 6184</lparam>
<lparam>Address:1829 6185</lparam>
<lparam>Address:1830 6192</lparam>
<lparam>Address:1831 6193</lparam>
<lparam>Address:1832 6194</lparam>
<lparam>Address:1833 6195</lparam>
<lparam>Address:1834 6196</lparam>
<lparam>Address:1835 6197</lparam>
<lparam>Address:1836 6198</lparam>
<lparam>Address:1837 6199</lparam>
<lparam>Address:1838 6200</lparam>
<lparam>Address:1839 6201</lparam>
<lparam>Address:1840 6208</lparam>
<lparam>Address:1841 6209</lparam>
<lparam>Address:1842 6210</lparam>
<lparam>Address:1843 6211</lparam>
<lparam>Address:1844 6212</lparam>
<lparam>Address:1845 6213</lparam>
<lparam>Address:1846 6214</lparam>
<lparam>Address:1847 6215</lparam>
<lparam>Address:1848 6216</lparam>
<lparam>Address:1849 6217</lparam>
<lparam>Address:1850 6224</lparam>
<lparam>Address:1851 6225</lparam>
<lparam>Address:1852 6226</lparam>
<lparam>Address:1853 6227</lparam>
<lparam>Address:1854 6228</lparam>
<lparam>Address:1855 6229</lparam>
<lparam>Address:1856 6230</lparam>
<lparam>Address:1857 6231</lparam>
<lparam>Address:1858 6232</lparam>
<lparam>Address:1859 6233</lparam>
<lparam>Address:1860 6240</lparam>
<lparam>Address:1861 6241</lparam>
<lparam>Address:1862 6242</lparam>
<lparam>Address:1863 6243</lparam>
<lparam>Address:1864 6244</lparam>
<lparam>Address:1865 6245</lparam>
<lparam>Address:1866 6246</lparam>
<lparam>Address:1867 6247</lparam>
<lparam>Address:1868 6248</lparam>
<lparam>Address:1869 6249</lparam>
<lparam>Address:1870 6256</lparam>
<lparam>Address:1871 6257</lparam>
<lparam>Address:1872 6258</lparam>
<lparam>Address:1873 6259</lparam>
<lparam>Address:1874 6260</lparam>
<lparam>Address:1875 6261</lparam>
<lparam>Address:1876 6262</lparam>
<lparam>Address:1877 6263</lparam>
<lparam>Address:1878 6264</lparam>
<lparam>Address:1879 6265</lparam>
<lparam>Address:1880 6272</lparam>
<lparam>Address:1881 6273</lparam>
<lparam>Address:1882 6274</lparam>
<lparam>Address:1883 6275</lparam>
<lparam>Address:1884 6276</lparam>
<lparam>Address:1885 6277</lparam>
<lparam>Address:1886 6278</lparam>
<lparam>Address:1887 6279</lparam>
<lparam>Address:1888 6280</lparam>
<lparam>Address:1889 6281</lparam>
<lparam>Address:1890 6288</lparam>
<lparam>Address:1891 6289</lparam>
<lparam>Address:1892 6290</lparam>
<lparam>Address:1893 6291</lparam>
<lparam>Address:1894 6292</lparam>
<lparam>Address:1895 6293</lparam>
<lparam>Address:1896 6294</lparam>
<lparam>Address:1897 6295</lparam>
<lparam>Address:1898 6296</lparam>
<lparam>Address:1899 6297</lparam>
<lparam>Address:1900 6400</lparam>
<lparam>Address:1901 6401</lparam>
<lparam>Address:1902 6402</lparam>
<lparam>Address:1903 6403</lparam>
<lparam>Address:1904 6404</lparam>
<lparam>Address:1905 6405</lparam>
<lparam>Address:1906 6406</lparam>
<lparam>Address:1907 6407</lparam>
<lparam>Address:1908 6408</lparam>
<lparam>Address:1909 6409</lparam>
<lparam>Address:1910 6416</lparam>
<lparam>Address:1911 6417</lparam>
<lparam>Address:1912 6418</lparam>
<lparam>Address:1913 6419</lparam>
<lparam>Address:1914 6420</lparam>
<lparam>Address:1915 6421</lparam>
<lparam>Address:1916 6422</lparam>
<lparam>Address:1917 6423</lparam>
<lparam>Address:1918 6424</lparam>
<lparam>Address:1919 6425</lparam>
<lparam>Address:1920 6432</lparam>
<lparam>Address:1921 6433</lparam>
<lparam>Address:1922 6434</lparam>
<lparam>Address:1923 6435</lparam>
<lparam>Address:1924 6436</lparam>
<lparam>Address:1925 6437</lparam>
<lparam>Address:1926 6438</lparam>
<lparam>Address:1927 6439</lparam>
<lparam>Address:1928 6440</lparam>
<lparam>Address:1929 6441</lparam>
<lparam>Address:1930 6448</lparam>
<lparam>Address:1931 6449</lparam>
<lparam>Address:1932 6450</lparam>
<lparam>Address:1933 6451</lparam>
<lparam>Address:1934 6452</lparam>
<lparam>Address:1935 6453</lparam>
<lparam>Address:1936 6454</lparam>
<lparam>Address:1937 6455</lparam>
<lparam>Address:1938 6456</lparam>
<lparam>Address:1939 6457</lparam>
<lparam>Address:1940 6464</lparam>
<lparam>Address:1941 6465</lparam>
<lparam>Address:1942 6466</lparam>
<lparam>Address:1943 6467</lparam>
<lparam>Address:1944 6468</lparam>
<lparam>Address:1945 6469</lparam>
<lparam>Address:1946 6470</lparam>
<lparam>Address:1947 6471</lparam>
<lparam>Address:1948 6472</lparam>
<lparam>Address:1949 6473</lparam>
<lparam>Address:1950 6480</lparam>
<lparam>Address:1951 6481</lparam>
<lparam>Address:1952 6482</lparam>
<lparam>Address:1953 6483</lparam>
<lparam>Address:1954 6484</lparam>
<lparam>Address:1955 6485</lparam>
<lparam>Address:1956 6486</lparam>
<lparam>Address:1957 6487</lparam>
<lparam>Address:1958 6488</lparam>
<lparam>Address:1959 6489</lparam>
<lparam>Address:1960 6496</lparam>
<lparam>Address:1961 6497</lparam>
<lparam>Address:1962 6498</lparam>
<lparam>Address:1963 6499</lparam>
<lparam>Address:1964 6500</lparam>
<lparam>Address:1965 6501</lparam>
<lparam>Address:1966 6502</lparam>
<lparam>Address:1967 6503</lparam>
<lparam>Address:1968 6504</lparam>
<lparam>Address:1969 6505</lparam>
<lparam>Address:1970 6512</lparam>
<lparam>Address:1971 6513</lparam>
<lparam>Address:1972 6514</lparam>
<lparam>Address:1973 6515</lparam>
<lparam>Address:1974 6516</lparam>
<lparam>Address:1975 6517</lparam>
<lparam>Address:1976 6518</lparam>
<lparam>Address:1977 6519</lparam>
<lparam>Address:1978 6520</lparam>
<lparam>Address:1979 6521</lparam>
<lparam>Address:1980 6528</lparam>
<lparam>Address:1981 6529</lparam>
<lparam>Address:1982 6530</lparam>
<lparam>Address:1983 6531</lparam>
<lparam>Address:1984 6532</lparam>
<lparam>Address:1985 6533</lparam>
<lparam>Address:1986 6534</lparam>
<lparam>Address:1987 6535</lparam>
<lparam>Address:1988 6536</lparam>
<lparam>Address:1989 6537</lparam>
<lparam>Address:1990 6544</lparam>
<lparam>Address:1991 6545</lparam>
<lparam>Address:1992 6546</lparam>
<lparam>Address:1993 6547</lparam>
<lparam>Address:1994 6548</lparam>
<lparam>Address:1995 6549</lparam>
<lparam>Address:1996 6550</lparam>
<lparam>Address:1997 6551</lparam>
<lparam>Address:1998 6552</lparam>
<lparam>Address:1999 6553</lparam>
<lparam>Address:2000 4096</lparam>
<lparam>Address:2001 8193</lparam>
<lparam>Address:2002 8194</lparam>
<lparam>Address:2003 8195</lparam>
<lparam>Address:2004 8196</lparam>
<lparam>Address:2005 8197</lparam>
<lparam>Address:2006 8198</lparam>
<lparam>Address:2007 8199</lparam>
<lparam>Address:2008 8200</lparam>
<lparam>Address:2009 8201</lparam>
<lparam>Address:2010 8208</lparam>
<lparam>Address:2011 8209</lparam>
<lparam>Address:2012 8210</lparam>
<lparam>Address:2013 8211</lparam>
<lparam>Address:2014 8212</lparam>
<lparam>Address:2015 8213</lparam>
<lparam>Address:2016 8214</lparam>
<lparam>Address:2017 8215</lparam>
<lparam>Address:2018 8216</lparam>
<lparam>Address:2019 8217</lparam>
<lparam>Address:2020 8224</lparam>
<lparam>Address:2021 8225</lparam>
<lparam>Address:2022 8226</lparam>
<lparam>Address:2023 8227</lparam>
<lparam>Address:2024 8228</lparam>
<lparam>Address:2025 8229</lparam>
<lparam>Address:2026 8230</lparam>
<lparam>Address:2027 8231</lparam>
<lparam>Address:2028 8232</lparam>
<lparam>Address:2029 8233</lparam>
<lparam>Address:2030 8240</lparam>
<lparam>Address:2031 8241</lparam>
<lparam>Address:2032 8242</lparam>
<lparam>Address:2033 8243</lparam>
<lparam>Address:2034 8244</lparam>
<lparam>Address:2035 8245</lparam>
<lparam>Address:2036 8246</lparam>
<lparam>Address:2037 8247</lparam>
<lparam>Address:2038 8248</lparam>
<lparam>Address:2039 8249</lparam>
<lparam>Address:2040 8256</lparam>
<lparam>Address:2041 8257</lparam>
<lparam>Address:2042 8258</lparam>
<lparam>Address:2043 8259</lparam>
<lparam>Address:2044 8260</lparam>
<lparam>Address:2045 8261</lparam>
<lparam>Address:2046 8262</lparam>
<lparam>Address:2047 8263</lparam>
<lparam>Address:2048 8264</lparam>
<lparam>Address:2049 8265</lparam>
<lparam>Address:2050 8272</lparam>
<lparam>Address:2051 8273</lparam>
<lparam>Address:2052 8274</lparam>
<lparam>Address:2053 8275</lparam>
<lparam>Address:2054 8276</lparam>
<lparam>Address:2055 8277</lparam>
<lparam>Address:2056 8278</lparam>
<lparam>Address:2057 8279</lparam>
<lparam>Address:2058 8280</lparam>
<lparam>Address:2059 8281</lparam>
<lparam>Address:2060 8288</lparam>
<lparam>Address:2061 8289</lparam>
<lparam>Address:2062 8290</lparam>
<lparam>Address:2063 8291</lparam>
<lparam>Address:2064 8292</lparam>
<lparam>Address:2065 8293</lparam>
<lparam>Address:2066 8294</lparam>
<lparam>Address:2067 8295</lparam>
<lparam>Address:2068 8296</lparam>
<lparam>Address:2069 8297</lparam>
<lparam>Address:2070 8304</lparam>
<lparam>Address:2071 8305</lparam>
<lparam>Address:2072 8306</lparam>
<lparam>Address:2073 8307</lparam>
<lparam>Address:2074 8308</lparam>
<lparam>Address:2075 8309</lparam>
<lparam>Address:2076 8310</lparam>
<lparam>Address:2077 8311</lparam>
<lparam>Address:2078 8312</lparam>
<lparam>Address:2079 8313</lparam>
<lparam>Address:2080 8320</lparam>
<lparam>Address:2081 8321</lparam>
<lparam>Address:2082 8322</lparam>
<lparam>Address:2083 8323</lparam>
<lparam>Address:2084 8324</lparam>
<lparam>Address:2085 8325</lparam>
<lparam>Address:2086 8326</lparam>
<lparam>Address:2087 8327</lparam>
<lparam>Address:2088 8328</lparam>
<lparam>Address:2089 8329</lparam>
<lparam>Address:2090 8336</lparam>
<lparam>Address:2091 8337</lparam>
<lparam>Address:2092 8338</lparam>
<lparam>Address:2093 8339</lparam>
<lparam>Address:2094 8340</lparam>
<lparam>Address:2095 8341</lparam>
<lparam>Address:2096 8342</lparam>
<lparam>Address:2097 8343</lparam>
<lparam>Address:2098 8344</lparam>
<lparam>Address:2099 8345</lparam>
<lparam>Address:2100 8448</lparam>
<lparam>Address:2101 8449</lparam>
<lparam>Address:2102 8450</lparam>
<lparam>Address:2103 8451</lparam>
<lparam>Address:2104 8452</lparam>
<lparam>Address:2105 8453</lparam>
<lparam>Address:2106 8454</lparam>
<lparam>Address:2107 8455</lparam>
<lparam>Address:2108 8456</lparam>
<lparam>Address:2109 8457</lparam>
<lparam>Address:2110 8464</lparam>
<lparam>Address:2111 8465</lparam>
<lparam>Address:2112 8466</lparam>
<lparam>Address:2113 8467</lparam>
<lparam>Address:2114 8468</lparam>
<lparam>Address:2115 8469</lparam>
<lparam>Address:2116 8470</lparam>
<lparam>Address:2117 8471</lparam>
<lparam>Address:2118 8472</lparam>
<lparam>Address:2119 8473</lparam>
<lparam>Address:2120 8480</lparam>
<lparam>Address:2121 8481</lparam>
<lparam>Address:2122 8482</lparam>
<lparam>Address:2123 8483</lparam>
<lparam>Address:2124 8484</lparam>
<lparam>Address:2125 8485</lparam>
<lparam>Address:2126 8486</lparam>
<lparam>Address:2127 8487</lparam>
<lparam>Address:2128 8488</lparam>
<lparam>Address:2129 8489</lparam>
<lparam>Address:2130 8496</lparam>
<lparam>Address:2131 8497</lparam>
<lparam>Address:2132 8498</lparam>
<lparam>Address:2133 8499</lparam>
<lparam>Address:2134 8500</lparam>
<lparam>Address:2135 8501</lparam>
<lparam>Address:2136 8502</lparam>
<lparam>Address:2137 8503</lparam>
<lparam>Address:2138 8504</lparam>
<lparam>Address:2139 8505</lparam>
<lparam>Address:2140 8512</lparam>
<lparam>Address:2141 8513</lparam>
<lparam>Address:2142 8514</lparam>
<lparam>Address:2143 8515</lparam>
<lparam>Address:2144 8516</lparam>
<lparam>Address:2145 8517</lparam>
<lparam>Address:2146 8518</lparam>
<lparam>Address:2147 8519</lparam>
<lparam>Address:2148 8520</lparam>
<lparam>Address:2149 8521</lparam>
<lparam>Address:2150 8528</lparam>
<lparam>Address:2151 8529</lparam>
<lparam>Address:2152 8530</lparam>
<lparam>Address:2153 8531</lparam>
<lparam>Address:2154 8532</lparam>
<lparam>Address:2155 8533</lparam>
<lparam>Address:2156 8534</lparam>
<lparam>Address:2157 8535</lparam>
<lparam>Address:2158 8536</lparam>
<lparam>Address:2159 8537</lparam>
<lparam>Address:2160 8544</lparam>
<lparam>Address:2161 8545</lparam>
<lparam>Address:2162 8546</lparam>
<lparam>Address:2163 8547</lparam>
<lparam>Address:2164 8548</lparam>
<lparam>Address:2165 8549</lparam>
<lparam>Address:2166 8550</lparam>
<lparam>Address:2167 8551</lparam>
<lparam>Address:2168 8552</lparam>
<lparam>Address:2169 8553</lparam>
<lparam>Address:2170 8560</lparam>
<lparam>Address:2171 8561</lparam>
<lparam>Address:2172 8562</lparam>
<lparam>Address:2173 8563</lparam>
<lparam>Address:2174 8564</lparam>
<lparam>Address:2175 8565</lparam>
<lparam>Address:2176 8566</lparam>
<lparam>Address:2177 8567</lparam>
<lparam>Address:2178 8568</lparam>
<lparam>Address:2179 8569</lparam>
<lparam>Address:2180 8576</lparam>
<lparam>Address:2181 8577</lparam>
<lparam>Address:2182 8578</lparam>
<lparam>Address:2183 8579</lparam>
<lparam>Address:2184 8580</lparam>
<lparam>Address:2185 8581</lparam>
<lparam>Address:2186 8582</lparam>
<lparam>Address:2187 8583</lparam>
<lparam>Address:2188 8584</lparam>
<lparam>Address:2189 8585</lparam>
<lparam>Address:2190 8592</lparam>
<lparam>Address:2191 8593</lparam>
<lparam>Address:2192 8594</lparam>
<lparam>Address:2193 8595</lparam>
<lparam>Address:2194 8596</lparam>
<lparam>Address:2195 8597</lparam>
<lparam>Address:2196 8598</lparam>
<lparam>Address:2197 8599</lparam>
<lparam>Address:2198 8600</lparam>
<lparam>Address:2199 8601</lparam>
<lparam>Address:2200 8704</lparam>
<lparam>Address:2201 8705</lparam>
<lparam>Address:2202 8706</lparam>
<lparam>Address:2203 8707</lparam>
<lparam>Address:2204 8708</lparam>
<lparam>Address:2205 8709</lparam>
<lparam>Address:2206 8710</lparam>
<lparam>Address:2207 8711</lparam>
<lparam>Address:2208 8712</lparam>
<lparam>Address:2209 8713</lparam>
<lparam>Address:2210 8720</lparam>
<lparam>Address:2211 8721</lparam>
<lparam>Address:2212 8722</lparam>
<lparam>Address:2213 8723</lparam>
<lparam>Address:2214 8724</lparam>
<lparam>Address:2215 8725</lparam>
<lparam>Address:2216 8726</lparam>
<lparam>Address:2217 8727</lparam>
<lparam>Address:2218 8728</lparam>
<lparam>Address:2219 8729</lparam>
<lparam>Address:2220 8736</lparam>
<lparam>Address:2221 8737</lparam>
<lparam>Address:2222 8738</lparam>
<lparam>Address:2223 8739</lparam>
<lparam>Address:2224 8740</lparam>
<lparam>Address:2225 8741</lparam>
<lparam>Address:2226 8742</lparam>
<lparam>Address:2227 8743</lparam>
<lparam>Address:2228 8744</lparam>
<lparam>Address:2229 8745</lparam>
<lparam>Address:2230 8752</lparam>
<lparam>Address:2231 8753</lparam>
<lparam>Address:2232 8754</lparam>
<lparam>Address:2233 8755</lparam>
<lparam>Address:2234 8756</lparam>
<lparam>Address:2235 8757</lparam>
<lparam>Address:2236 8758</lparam>
<lparam>Address:2237 8759</lparam>
<lparam>Address:2238 8760</lparam>
<lparam>Address:2239 8761</lparam>
<lparam>Address:2240 8768</lparam>
<lparam>Address:2241 8769</lparam>
<lparam>Address:2242 8770</lparam>
<lparam>Address:2243 8771</lparam>
<lparam>Address:2244 8772</lparam>
<lparam>Address:2245 8773</lparam>
<lparam>Address:2246 8774</lparam>
<lparam>Address:2247 8775</lparam>
<lparam>Address:2248 8776</lparam>
<lparam>Address:2249 8777</lparam>
<lparam>Address:2250 8784</lparam>
<lparam>Address:2251 8785</lparam>
<lparam>Address:2252 8786</lparam>
<lparam>Address:2253 8787</lparam>
<lparam>Address:2254 8788</lparam>
<lparam>Address:2255 8789</lparam>
<lparam>Address:2256 8790</lparam>
<lparam>Address:2257 8791</lparam>
<lparam>Address:2258 8792</lparam>
<lparam>Address:2259 8793</lparam>
<lparam>Address:2260 8800</lparam>
<lparam>Address:2261 8801</lparam>
<lparam>Address:2262 8802</lparam>
<lparam>Address:2263 8803</lparam>
<lparam>Address:2264 8804</lparam>
<lparam>Address:2265 8805</lparam>
<lparam>Address:2266 8806</lparam>
<lparam>Address:2267 8807</lparam>
<lparam>Address:2268 8808</lparam>
<lparam>Address:2269 8809</lparam>
<lparam>Address:2270 8816</lparam>
<lparam>Address:2271 8817</lparam>
<lparam>Address:2272 8818</lparam>
<lparam>Address:2273 8819</lparam>
<lparam>Address:2274 8820</lparam>
<lparam>Address:2275 8821</lparam>
<lparam>Address:2276 8822</lparam>
<lparam>Address:2277 8823</lparam>
<lparam>Address:2278 8824</lparam>
<lparam>Address:2279 8825</lparam>
<lparam>Address:2280 8832</lparam>
<lparam>Address:2281 8833</lparam>
<lparam>Address:2282 8834</lparam>
<lparam>Address:2283 8835</lparam>
<lparam>Address:2284 8836</lparam>
<lparam>Address:2285 8837</lparam>
<lparam>Address:2286 8838</lparam>
<lparam>Address:2287 8839</lparam>
<lparam>Address:2288 8840</lparam>
<lparam>Address:2289 8841</lparam>
<lparam>Address:2290 8848</lparam>
<lparam>Address:2291 8849</lparam>
<lparam>Address:2292 8850</lparam>
<lparam>Address:2293 8851</lparam>
<lparam>Address:2294 8852</lparam>
<lparam>Address:2295 8853</lparam>
<lparam>Address:2296 8854</lparam>
<lparam>Address:2297 8855</lparam>
<lparam>Address:2298 8856</lparam>
<lparam>Address:2299 8857</lparam>
<lparam>Address:2300 8960</lparam>
<lparam>Address:2301 8961</lparam>
<lparam>Address:2302 8962</lparam>
<lparam>Address:2303 8963</lparam>
<lparam>Address:2304 8964</lparam>
<lparam>Address:2305 8965</lparam>
<lparam>Address:2306 8966</lparam>
<lparam>Address:2307 8967</lparam>
<lparam>Address:2308 8968</lparam>
<lparam>Address:2309 8969</lparam>
<lparam>Address:2310 8976</lparam>
<lparam>Address:2311 8977</lparam>
<lparam>Address:2312 8978</lparam>
<lparam>Address:2313 8979</lparam>
<lparam>Address:2314 8980</lparam>
<lparam>Address:2315 8981</lparam>
<lparam>Address:2316 8982</lparam>
<lparam>Address:2317 8983</lparam>
<lparam>Address:2318 8984</lparam>
<lparam>Address:2319 8985</lparam>
<lparam>Address:2320 8992</lparam>
<lparam>Address:2321 8993</lparam>
<lparam>Address:2322 8994</lparam>
<lparam>Address:2323 8995</lparam>
<lparam>Address:2324 8996</lparam>
<lparam>Address:2325 8997</lparam>
<lparam>Address:2326 8998</lparam>
<lparam>Address:2327 8999</lparam>
<lparam>Address:2328 9000</lparam>
<lparam>Address:2329 9001</lparam>
<lparam>Address:2330 9008</lparam>
<lparam>Address:2331 9009</lparam>
<lparam>Address:2332 9010</lparam>
<lparam>Address:2333 9011</lparam>
<lparam>Address:2334 9012</lparam>
<lparam>Address:2335 9013</lparam>
<lparam>Address:2336 9014</lparam>
<lparam>Address:2337 9015</lparam>
<lparam>Address:2338 9016</lparam>
<lparam>Address:2339 9017</lparam>
<lparam>Address:2340 9024</lparam>
<lparam>Address:2341 9025</lparam>
<lparam>Address:2342 9026</lparam>
<lparam>Address:2343 9027</lparam>
<lparam>Address:2344 9028</lparam>
<lparam>Address:2345 9029</lparam>
<lparam>Address:2346 9030</lparam>
<lparam>Address:2347 9031</lparam>
<lparam>Address:2348 9032</lparam>
<lparam>Address:2349 9033</lparam>
<lparam>Address:2350 9040</lparam>
<lparam>Address:2351 9041</lparam>
<lparam>Address:2352 9042</lparam>
<lparam>Address:2353 9043</lparam>
<lparam>Address:2354 9044</lparam>
<lparam>Address:2355 9045</lparam>
<lparam>Address:2356 9046</lparam>
<lparam>Address:2357 9047</lparam>
<lparam>Address:2358 9048</lparam>
<lparam>Address:2359 9049</lparam>
<lparam>Address:2360 9056</lparam>
<lparam>Address:2361 9057</lparam>
<lparam>Address:2362 9058</lparam>
<lparam>Address:2363 9059</lparam>
<lparam>Address:2364 9060</lparam>
<lparam>Address:2365 9061</lparam>
<lparam>Address:2366 9062</lparam>
<lparam>Address:2367 9063</lparam>
<lparam>Address:2368 9064</lparam>
<lparam>Address:2369 9065</lparam>
<lparam>Address:2370 9072</lparam>
<lparam>Address:2371 9073</lparam>
<lparam>Address:2372 9074</lparam>
<lparam>Address:2373 9075</lparam>
<lparam>Address:2374 9076</lparam>
<lparam>Address:2375 9077</lparam>
<lparam>Address:2376 9078</lparam>
<lparam>Address:2377 9079</lparam>
<lparam>Address:2378 9080</lparam>
<lparam>Address:2379 9081</lparam>
<lparam>Address:2380 9088</lparam>
<lparam>Address:2381 9089</lparam>
<lparam>Address:2382 9090</lparam>
<lparam>Address:2383 9091</lparam>
<lparam>Address:2384 9092</lparam>
<lparam>Address:2385 9093</lparam>
<lparam>Address:2386 9094</lparam>
<lparam>Address:2387 9095</lparam>
<lparam>Address:2388 9096</lparam>
<lparam>Address:2389 9097</lparam>
<lparam>Address:2390 9104</lparam>
<lparam>Address:2391 9105</lparam>
<lparam>Address:2392 9106</lparam>
<lparam>Address:2393 9107</lparam>
<lparam>Address:2394 9108</lparam>
<lparam>Address:2395 9109</lparam>
<lparam>Address:2396 9110</lparam>
<lparam>Address:2397 9111</lparam>
<lparam>Address:2398 9112</lparam>
<lparam>Address:2399 9113</lparam>
<lparam>Address:2400 9216</lparam>
<lparam>Address:2401 9217</lparam>
<lparam>Address:2402 9218</lparam>
<lparam>Address:2403 9219</lparam>
<lparam>Address:2404 9220</lparam>
<lparam>Address:2405 9221</lparam>
<lparam>Address:2406 9222</lparam>
<lparam>Address:2407 9223</lparam>
<lparam>Address:2408 9224</lparam>
<lparam>Address:2409 9225</lparam>
<lparam>Address:2410 9232</lparam>
<lparam>Address:2411 9233</lparam>
<lparam>Address:2412 9234</lparam>
<lparam>Address:2413 9235</lparam>
<lparam>Address:2414 9236</lparam>
<lparam>Address:2415 9237</lparam>
<lparam>Address:2416 9238</lparam>
<lparam>Address:2417 9239</lparam>
<lparam>Address:2418 9240</lparam>
<lparam>Address:2419 9241</lparam>
<lparam>Address:2420 9248</lparam>
<lparam>Address:2421 9249</lparam>
<lparam>Address:2422 9250</lparam>
<lparam>Address:2423 9251</lparam>
<lparam>Address:2424 9252</lparam>
<lparam>Address:2425 9253</lparam>
<lparam>Address:2426 9254</lparam>
<lparam>Address:2427 9255</lparam>
<lparam>Address:2428 9256</lparam>
<lparam>Address:2429 9257</lparam>
<lparam>Address:2430 9264</lparam>
<lparam>Address:2431 9265</lparam>
<lparam>Address:2432 9266</lparam>
<lparam>Address:2433 9267</lparam>
<lparam>Address:2434 9268</lparam>
<lparam>Address:2435 9269</lparam>
<lparam>Address:2436 9270</lparam>
<lparam>Address:2437 9271</lparam>
<lparam>Address:2438 9272</lparam>
<lparam>Address:2439 9273</lparam>
<lparam>Address:2440 9280</lparam>
<lparam>Address:2441 9281</lparam>
<lparam>Address:2442 9282</lparam>
<lparam>Address:2443 9283</lparam>
<lparam>Address:2444 9284</lparam>
<lparam>Address:2445 9285</lparam>
<lparam>Address:2446 9286</lparam>
<lparam>Address:2447 9287</lparam>
<lparam>Address:2448 9288</lparam>
<lparam>Address:2449 9289</lparam>
<lparam>Address:2450 9296</lparam>
<lparam>Address:2451 9297</lparam>
<lparam>Address:2452 9298</lparam>
<lparam>Address:2453 9299</lparam>
<lparam>Address:2454 9300</lparam>
<lparam>Address:2455 9301</lparam>
<lparam>Address:2456 9302</lparam>
<lparam>Address:2457 9303</lparam>
<lparam>Address:2458 9304</lparam>
<lparam>Address:2459 9305</lparam>
<lparam>Address:2460 9312</lparam>
<lparam>Address:2461 9313</lparam>
<lparam>Address:2462 9314</lparam>
<lparam>Address:2463 9315</lparam>
<lparam>Address:2464 9316</lparam>
<lparam>Address:2465 9317</lparam>
<lparam>Address:2466 9318</lparam>
<lparam>Address:2467 9319</lparam>
<lparam>Address:2468 9320</lparam>
<lparam>Address:2469 9321</lparam>
<lparam>Address:2470 9328</lparam>
<lparam>Address:2471 9329</lparam>
<lparam>Address:2472 9330</lparam>
<lparam>Address:2473 9331</lparam>
<lparam>Address:2474 9332</lparam>
<lparam>Address:2475 9333</lparam>
<lparam>Address:2476 9334</lparam>
<lparam>Address:2477 9335</lparam>
<lparam>Address:2478 9336</lparam>
<lparam>Address:2479 9337</lparam>
<lparam>Address:2480 9344</lparam>
<lparam>Address:2481 9345</lparam>
<lparam>Address:2482 9346</lparam>
<lparam>Address:2483 9347</lparam>
<lparam>Address:2484 9348</lparam>
<lparam>Address:2485 9349</lparam>
<lparam>Address:2486 9350</lparam>
<lparam>Address:2487 9351</lparam>
<lparam>Address:2488 9352</lparam>
<lparam>Address:2489 9353</lparam>
<lparam>Address:2490 9360</lparam>
<lparam>Address:2491 9361</lparam>
<lparam>Address:2492 9362</lparam>
<lparam>Address:2493 9363</lparam>
<lparam>Address:2494 9364</lparam>
<lparam>Address:2495 9365</lparam>
<lparam>Address:2496 9366</lparam>
<lparam>Address:2497 9367</lparam>
<lparam>Address:2498 9368</lparam>
<lparam>Address:2499 9369</lparam>
<lparam>Address:2500 9472</lparam>
<lparam>Address:2501 9473</lparam>
<lparam>Address:2502 9474</lparam>
<lparam>Address:2503 9475</lparam>
<lparam>Address:2504 9476</lparam>
<lparam>Address:2505 9477</lparam>
<lparam>Address:2506 9478</lparam>
<lparam>Address:2507 9479</lparam>
<lparam>Address:2508 9480</lparam>
<lparam>Address:2509 9481</lparam>
<lparam>Address:2510 9488</lparam>
<lparam>Address:2511 9489</lparam>
<lparam>Address:2512 9490</lparam>
<lparam>Address:2513 9491</lparam>
<lparam>Address:2514 9492</lparam>
<lparam>Address:2515 9493</lparam>
<lparam>Address:2516 9494</lparam>
<lparam>Address:2517 9495</lparam>
<lparam>Address:2518 9496</lparam>
<lparam>Address:2519 9497</lparam>
<lparam>Address:2520 9504</lparam>
<lparam>Address:2521 9505</lparam>
<lparam>Address:2522 9506</lparam>
<lparam>Address:2523 9507</lparam>
<lparam>Address:2524 9508</lparam>
<lparam>Address:2525 9509</lparam>
<lparam>Address:2526 9510</lparam>
<lparam>Address:2527 9511</lparam>
<lparam>Address:2528 9512</lparam>
<lparam>Address:2529 9513</lparam>
<lparam>Address:2530 9520</lparam>
<lparam>Address:2531 9521</lparam>
<lparam>Address:2532 9522</lparam>
<lparam>Address:2533 9523</lparam>
<lparam>Address:2534 9524</lparam>
<lparam>Address:2535 9525</lparam>
<lparam>Address:2536 9526</lparam>
<lparam>Address:2537 9527</lparam>
<lparam>Address:2538 9528</lparam>
<lparam>Address:2539 9529</lparam>
<lparam>Address:2540 9536</lparam>
<lparam>Address:2541 9537</lparam>
<lparam>Address:2542 9538</lparam>
<lparam>Address:2543 9539</lparam>
<lparam>Address:2544 9540</lparam>
<lparam>Address:2545 9541</lparam>
<lparam>Address:2546 9542</lparam>
<lparam>Address:2547 9543</lparam>
<lparam>Address:2548 9544</lparam>
<lparam>Address:2549 9545</lparam>
<lparam>Address:2550 9552</lparam>
<lparam>Address:2551 9553</lparam>
<lparam>Address:2552 9554</lparam>
<lparam>Address:2553 9555</lparam>
<lparam>Address:2554 9556</lparam>
<lparam>Address:2555 9557</lparam>
<lparam>Address:2556 9558</lparam>
<lparam>Address:2557 9559</lparam>
<lparam>Address:2558 9560</lparam>
<lparam>Address:2559 9561</lparam>
<lparam>Address:2560 9568</lparam>
<lparam>Address:2561 9569</lparam>
<lparam>Address:2562 9570</lparam>
<lparam>Address:2563 9571</lparam>
<lparam>Address:2564 9572</lparam>
<lparam>Address:2565 9573</lparam>
<lparam>Address:2566 9574</lparam>
<lparam>Address:2567 9575</lparam>
<lparam>Address:2568 9576</lparam>
<lparam>Address:2569 9577</lparam>
<lparam>Address:2570 9584</lparam>
<lparam>Address:2571 9585</lparam>
<lparam>Address:2572 9586</lparam>
<lparam>Address:2573 9587</lparam>
<lparam>Address:2574 9588</lparam>
<lparam>Address:2575 9589</lparam>
<lparam>Address:2576 9590</lparam>
<lparam>Address:2577 9591</lparam>
<lparam>Address:2578 9592</lparam>
<lparam>Address:2579 9593</lparam>
<lparam>Address:2580 9600</lparam>
<lparam>Address:2581 9601</lparam>
<lparam>Address:2582 9602</lparam>
<lparam>Address:2583 9603</lparam>
<lparam>Address:2584 9604</lparam>
<lparam>Address:2585 9605</lparam>
<lparam>Address:2586 9606</lparam>
<lparam>Address:2587 9607</lparam>
<lparam>Address:2588 9608</lparam>
<lparam>Address:2589 9609</lparam>
<lparam>Address:2590 9616</lparam>
<lparam>Address:2591 9617</lparam>
<lparam>Address:2592 9618</lparam>
<lparam>Address:2593 9619</lparam>
<lparam>Address:2594 9620</lparam>
<lparam>Address:2595 9621</lparam>
<lparam>Address:2596 9622</lparam>
<lparam>Address:2597 9623</lparam>
<lparam>Address:2598 9624</lparam>
<lparam>Address:2599 9625</lparam>
<lparam>Address:2600 9728</lparam>
<lparam>Address:2601 9729</lparam>
<lparam>Address:2602 9730</lparam>
<lparam>Address:2603 9731</lparam>
<lparam>Address:2604 9732</lparam>
<lparam>Address:2605 9733</lparam>
<lparam>Address:2606 9734</lparam>
<lparam>Address:2607 9735</lparam>
<lparam>Address:2608 9736</lparam>
<lparam>Address:2609 9737</lparam>
<lparam>Address:2610 9744</lparam>
<lparam>Address:2611 9745</lparam>
<lparam>Address:2612 9746</lparam>
<lparam>Address:2613 9747</lparam>
<lparam>Address:2614 9748</lparam>
<lparam>Address:2615 9749</lparam>
<lparam>Address:2616 9750</lparam>
<lparam>Address:2617 9751</lparam>
<lparam>Address:2618 9752</lparam>
<lparam>Address:2619 9753</lparam>
<lparam>Address:2620 9760</lparam>
<lparam>Address:2621 9761</lparam>
<lparam>Address:2622 9762</lparam>
<lparam>Address:2623 9763</lparam>
<lparam>Address:2624 9764</lparam>
<lparam>Address:2625 9765</lparam>
<lparam>Address:2626 9766</lparam>
<lparam>Address:2627 9767</lparam>
<lparam>Address:2628 9768</lparam>
<lparam>Address:2629 9769</lparam>
<lparam>Address:2630 9776</lparam>
<lparam>Address:2631 9777</lparam>
<lparam>Address:2632 9778</lparam>
<lparam>Address:2633 9779</lparam>
<lparam>Address:2634 9780</lparam>
<lparam>Address:2635 9781</lparam>
<lparam>Address:2636 9782</lparam>
<lparam>Address:2637 9783</lparam>
<lparam>Address:2638 9784</lparam>
<lparam>Address:2639 9785</lparam>
<lparam>Address:2640 9792</lparam>
<lparam>Address:2641 9793</lparam>
<lparam>Address:2642 9794</lparam>
<lparam>Address:2643 9795</lparam>
<lparam>Address:2644 9796</lparam>
<lparam>Address:2645 9797</lparam>
<lparam>Address:2646 9798</lparam>
<lparam>Address:2647 9799</lparam>
<lparam>Address:2648 9800</lparam>
<lparam>Address:2649 9801</lparam>
<lparam>Address:2650 9808</lparam>
<lparam>Address:2651 9809</lparam>
<lparam>Address:2652 9810</lparam>
<lparam>Address:2653 9811</lparam>
<lparam>Address:2654 9812</lparam>
<lparam>Address:2655 9813</lparam>
<lparam>Address:2656 9814</lparam>
<lparam>Address:2657 9815</lparam>
<lparam>Address:2658 9816</lparam>
<lparam>Address:2659 9817</lparam>
<lparam>Address:2660 9824</lparam>
<lparam>Address:2661 9825</lparam>
<lparam>Address:2662 9826</lparam>
<lparam>Address:2663 9827</lparam>
<lparam>Address:2664 9828</lparam>
<lparam>Address:2665 9829</lparam>
<lparam>Address:2666 9830</lparam>
<lparam>Address:2667 9831</lparam>
<lparam>Address:2668 9832</lparam>
<lparam>Address:2669 9833</lparam>
<lparam>Address:2670 9840</lparam>
<lparam>Address:2671 9841</lparam>
<lparam>Address:2672 9842</lparam>
<lparam>Address:2673 9843</lparam>
<lparam>Address:2674 9844</lparam>
<lparam>Address:2675 9845</lparam>
<lparam>Address:2676 9846</lparam>
<lparam>Address:2677 9847</lparam>
<lparam>Address:2678 9848</lparam>
<lparam>Address:2679 9849</lparam>
<lparam>Address:2680 9856</lparam>
<lparam>Address:2681 9857</lparam>
<lparam>Address:2682 9858</lparam>
<lparam>Address:2683 9859</lparam>
<lparam>Address:2684 9860</lparam>
<lparam>Address:2685 9861</lparam>
<lparam>Address:2686 9862</lparam>
<lparam>Address:2687 9863</lparam>
<lparam>Address:2688 9864</lparam>
<lparam>Address:2689 9865</lparam>
<lparam>Address:2690 9872</lparam>
<lparam>Address:2691 9873</lparam>
<lparam>Address:2692 9874</lparam>
<lparam>Address:2693 9875</lparam>
<lparam>Address:2694 9876</lparam>
<lparam>Address:2695 9877</lparam>
<lparam>Address:2696 9878</lparam>
<lparam>Address:2697 9879</lparam>
<lparam>Address:2698 9880</lparam>
<lparam>Address:2699 9881</lparam>
<lparam>Address:2700 9984</lparam>
<lparam>Address:2701 9985</lparam>
<lparam>Address:2702 9986</lparam>
<lparam>Address:2703 9987</lparam>
<lparam>Address:2704 9988</lparam>
<lparam>Address:2705 9989</lparam>
<lparam>Address:2706 9990</lparam>
<lparam>Address:2707 9991</lparam>
<lparam>Address:2708 9992</lparam>
<lparam>Address:2709 9993</lparam>
<lparam>Address:2710 10000</lparam>
<lparam>Address:2711 10001</lparam>
<lparam>Address:2712 10002</lparam>
<lparam>Address:2713 10003</lparam>
<lparam>Address:2714 10004</lparam>
<lparam>Address:2715 10005</lparam>
<lparam>Address:2716 10006</lparam>
<lparam>Address:2717 10007</lparam>
<lparam>Address:2718 10008</lparam>
<lparam>Address:2719 10009</lparam>
<lparam>Address:2720 10016</lparam>
<lparam>Address:2721 10017</lparam>
<lparam>Address:2722 10018</lparam>
<lparam>Address:2723 10019</lparam>
<lparam>Address:2724 10020</lparam>
<lparam>Address:2725 10021</lparam>
<lparam>Address:2726 10022</lparam>
<lparam>Address:2727 10023</lparam>
<lparam>Address:2728 10024</lparam>
<lparam>Address:2729 10025</lparam>
<lparam>Address:2730 10032</lparam>
<lparam>Address:2731 10033</lparam>
<lparam>Address:2732 10034</lparam>
<lparam>Address:2733 10035</lparam>
<lparam>Address:2734 10036</lparam>
<lparam>Address:2735 10037</lparam>
<lparam>Address:2736 10038</lparam>
<lparam>Address:2737 10039</lparam>
<lparam>Address:2738 10040</lparam>
<lparam>Address:2739 10041</lparam>
<lparam>Address:2740 10048</lparam>
<lparam>Address:2741 10049</lparam>
<lparam>Address:2742 10050</lparam>
<lparam>Address:2743 10051</lparam>
<lparam>Address:2744 10052</lparam>
<lparam>Address:2745 10053</lparam>
<lparam>Address:2746 10054</lparam>
<lparam>Address:2747 10055</lparam>
<lparam>Address:2748 10056</lparam>
<lparam>Address:2749 10057</lparam>
<lparam>Address:2750 10064</lparam>
<lparam>Address:2751 10065</lparam>
<lparam>Address:2752 10066</lparam>
<lparam>Address:2753 10067</lparam>
<lparam>Address:2754 10068</lparam>
<lparam>Address:2755 10069</lparam>
<lparam>Address:2756 10070</lparam>
<lparam>Address:2757 10071</lparam>
<lparam>Address:2758 10072</lparam>
<lparam>Address:2759 10073</lparam>
<lparam>Address:2760 10080</lparam>
<lparam>Address:2761 10081</lparam>
<lparam>Address:2762 10082</lparam>
<lparam>Address:2763 10083</lparam>
<lparam>Address:2764 10084</lparam>
<lparam>Address:2765 10085</lparam>
<lparam>Address:2766 10086</lparam>
<lparam>Address:2767 10087</lparam>
<lparam>Address:2768 10088</lparam>
<lparam>Address:2769 10089</lparam>
<lparam>Address:2770 10096</lparam>
<lparam>Address:2771 10097</lparam>
<lparam>Address:2772 10098</lparam>
<lparam>Address:2773 10099</lparam>
<lparam>Address:2774 10100</lparam>
<lparam>Address:2775 10101</lparam>
<lparam>Address:2776 10102</lparam>
<lparam>Address:2777 10103</lparam>
<lparam>Address:2778 10104</lparam>
<lparam>Address:2779 10105</lparam>
<lparam>Address:2780 10112</lparam>
<lparam>Address:2781 10113</lparam>
<lparam>Address:2782 10114</lparam>
<lparam>Address:2783 10115</lparam>
<lparam>Address:2784 10116</lparam>
<lparam>Address:2785 10117</lparam>
<lparam>Address:2786 10118</lparam>
<lparam>Address:2787 10119</lparam>
<lparam>Address:2788 10120</lparam>
<lparam>Address:2789 10121</lparam>
<lparam>Address:2790 10128</lparam>
<lparam>Address:2791 10129</lparam>
<lparam>Address:2792 10130</lparam>
<lparam>Address:2793 10131</lparam>
<lparam>Address:2794 10132</lparam>
<lparam>Address:2795 10133</lparam>
<lparam>Address:2796 10134</lparam>
<lparam>Address:2797 10135</lparam>
<lparam>Address:2798 10136</lparam>
<lparam>Address:2799 10137</lparam>
<lparam>Address:2800 10240</lparam>
<lparam>Address:2801 10241</lparam>
<lparam>Address:2802 10242</lparam>
<lparam>Address:2803 10243</lparam>
<lparam>Address:2804 10244</lparam>
<lparam>Address:2805 10245</lparam>
<lparam>Address:2806 10246</lparam>
<lparam>Address:2807 10247</lparam>
<lparam>Address:2808 10248</lparam>
<lparam>Address:2809 10249</lparam>
<lparam>Address:2810 10256</lparam>
<lparam>Address:2811 10257</lparam>
<lparam>Address:2812 10258</lparam>
<lparam>Address:2813 10259</lparam>
<lparam>Address:2814 10260</lparam>
<lparam>Address:2815 10261</lparam>
<lparam>Address:2816 10262</lparam>
<lparam>Address:2817 10263</lparam>
<lparam>Address:2818 10264</lparam>
<lparam>Address:2819 10265</lparam>
<lparam>Address:2820 10272</lparam>
<lparam>Address:2821 10273</lparam>
<lparam>Address:2822 10274</lparam>
<lparam>Address:2823 10275</lparam>
<lparam>Address:2824 10276</lparam>
<lparam>Address:2825 10277</lparam>
<lparam>Address:2826 10278</lparam>
<lparam>Address:2827 10279</lparam>
<lparam>Address:2828 10280</lparam>
<lparam>Address:2829 10281</lparam>
<lparam>Address:2830 10288</lparam>
<lparam>Address:2831 10289</lparam>
<lparam>Address:2832 10290</lparam>
<lparam>Address:2833 10291</lparam>
<lparam>Address:2834 10292</lparam>
<lparam>Address:2835 10293</lparam>
<lparam>Address:2836 10294</lparam>
<lparam>Address:2837 10295</lparam>
<lparam>Address:2838 10296</lparam>
<lparam>Address:2839 10297</lparam>
<lparam>Address:2840 10304</lparam>
<lparam>Address:2841 10305</lparam>
<lparam>Address:2842 10306</lparam>
<lparam>Address:2843 10307</lparam>
<lparam>Address:2844 10308</lparam>
<lparam>Address:2845 10309</lparam>
<lparam>Address:2846 10310</lparam>
<lparam>Address:2847 10311</lparam>
<lparam>Address:2848 10312</lparam>
<lparam>Address:2849 10313</lparam>
<lparam>Address:2850 10320</lparam>
<lparam>Address:2851 10321</lparam>
<lparam>Address:2852 10322</lparam>
<lparam>Address:2853 10323</lparam>
<lparam>Address:2854 10324</lparam>
<lparam>Address:2855 10325</lparam>
<lparam>Address:2856 10326</lparam>
<lparam>Address:2857 10327</lparam>
<lparam>Address:2858 10328</lparam>
<lparam>Address:2859 10329</lparam>
<lparam>Address:2860 10336</lparam>
<lparam>Address:2861 10337</lparam>
<lparam>Address:2862 10338</lparam>
<lparam>Address:2863 10339</lparam>
<lparam>Address:2864 10340</lparam>
<lparam>Address:2865 10341</lparam>
<lparam>Address:2866 10342</lparam>
<lparam>Address:2867 10343</lparam>
<lparam>Address:2868 10344</lparam>
<lparam>Address:2869 10345</lparam>
<lparam>Address:2870 10352</lparam>
<lparam>Address:2871 10353</lparam>
<lparam>Address:2872 10354</lparam>
<lparam>Address:2873 10355</lparam>
<lparam>Address:2874 10356</lparam>
<lparam>Address:2875 10357</lparam>
<lparam>Address:2876 10358</lparam>
<lparam>Address:2877 10359</lparam>
<lparam>Address:2878 10360</lparam>
<lparam>Address:2879 10361</lparam>
<lparam>Address:2880 10368</lparam>
<lparam>Address:2881 10369</lparam>
<lparam>Address:2882 10370</lparam>
<lparam>Address:2883 10371</lparam>
<lparam>Address:2884 10372</lparam>
<lparam>Address:2885 10373</lparam>
<lparam>Address:2886 10374</lparam>
<lparam>Address:2887 10375</lparam>
<lparam>Address:2888 10376</lparam>
<lparam>Address:2889 10377</lparam>
<lparam>Address:2890 10384</lparam>
<lparam>Address:2891 10385</lparam>
<lparam>Address:2892 10386</lparam>
<lparam>Address:2893 10387</lparam>
<lparam>Address:2894 10388</lparam>
<lparam>Address:2895 10389</lparam>
<lparam>Address:2896 10390</lparam>
<lparam>Address:2897 10391</lparam>
<lparam>Address:2898 10392</lparam>
<lparam>Address:2899 10393</lparam>
<lparam>Address:2900 10496</lparam>
<lparam>Address:2901 10497</lparam>
<lparam>Address:2902 10498</lparam>
<lparam>Address:2903 10499</lparam>
<lparam>Address:2904 10500</lparam>
<lparam>Address:2905 10501</lparam>
<lparam>Address:2906 10502</lparam>
<lparam>Address:2907 10503</lparam>
<lparam>Address:2908 10504</lparam>
<lparam>Address:2909 10505</lparam>
<lparam>Address:2910 10512</lparam>
<lparam>Address:2911 10513</lparam>
<lparam>Address:2912 10514</lparam>
<lparam>Address:2913 10515</lparam>
<lparam>Address:2914 10516</lparam>
<lparam>Address:2915 10517</lparam>
<lparam>Address:2916 10518</lparam>
<lparam>Address:2917 10519</lparam>
<lparam>Address:2918 10520</lparam>
<lparam>Address:2919 10521</lparam>
<lparam>Address:2920 10528</lparam>
<lparam>Address:2921 10529</lparam>
<lparam>Address:2922 10530</lparam>
<lparam>Address:2923 10531</lparam>
<lparam>Address:2924 10532</lparam>
<lparam>Address:2925 10533</lparam>
<lparam>Address:2926 10534</lparam>
<lparam>Address:2927 10535</lparam>
<lparam>Address:2928 10536</lparam>
<lparam>Address:2929 10537</lparam>
<lparam>Address:2930 10544</lparam>
<lparam>Address:2931 10545</lparam>
<lparam>Address:2932 10546</lparam>
<lparam>Address:2933 10547</lparam>
<lparam>Address:2934 10548</lparam>
<lparam>Address:2935 10549</lparam>
<lparam>Address:2936 10550</lparam>
<lparam>Address:2937 10551</lparam>
<lparam>Address:2938 10552</lparam>
<lparam>Address:2939 10553</lparam>
<lparam>Address:2940 10560</lparam>
<lparam>Address:2941 10561</lparam>
<lparam>Address:2942 10562</lparam>
<lparam>Address:2943 10563</lparam>
<lparam>Address:2944 10564</lparam>
<lparam>Address:2945 10565</lparam>
<lparam>Address:2946 10566</lparam>
<lparam>Address:2947 10567</lparam>
<lparam>Address:2948 10568</lparam>
<lparam>Address:2949 10569</lparam>
<lparam>Address:2950 10576</lparam>
<lparam>Address:2951 10577</lparam>
<lparam>Address:2952 10578</lparam>
<lparam>Address:2953 10579</lparam>
<lparam>Address:2954 10580</lparam>
<lparam>Address:2955 10581</lparam>
<lparam>Address:2956 10582</lparam>
<lparam>Address:2957 10583</lparam>
<lparam>Address:2958 10584</lparam>
<lparam>Address:2959 10585</lparam>
<lparam>Address:2960 10592</lparam>
<lparam>Address:2961 10593</lparam>
<lparam>Address:2962 10594</lparam>
<lparam>Address:2963 10595</lparam>
<lparam>Address:2964 10596</lparam>
<lparam>Address:2965 10597</lparam>
<lparam>Address:2966 10598</lparam>
<lparam>Address:2967 10599</lparam>
<lparam>Address:2968 10600</lparam>
<lparam>Address:2969 10601</lparam>
<lparam>Address:2970 10608</lparam>
<lparam>Address:2971 10609</lparam>
<lparam>Address:2972 10610</lparam>
<lparam>Address:2973 10611</lparam>
<lparam>Address:2974 10612</lparam>
<lparam>Address:2975 10613</lparam>
<lparam>Address:2976 10614</lparam>
<lparam>Address:2977 10615</lparam>
<lparam>Address:2978 10616</lparam>
<lparam>Address:2979 10617</lparam>
<lparam>Address:2980 10624</lparam>
<lparam>Address:2981 10625</lparam>
<lparam>Address:2982 10626</lparam>
<lparam>Address:2983 10627</lparam>
<lparam>Address:2984 10628</lparam>
<lparam>Address:2985 10629</lparam>
<lparam>Address:2986 10630</lparam>
<lparam>Address:2987 10631</lparam>
<lparam>Address:2988 10632</lparam>
<lparam>Address:2989 10633</lparam>
<lparam>Address:2990 10640</lparam>
<lparam>Address:2991 10641</lparam>
<lparam>Address:2992 10642</lparam>
<lparam>Address:2993 10643</lparam>
<lparam>Address:2994 10644</lparam>
<lparam>Address:2995 10645</lparam>
<lparam>Address:2996 10646</lparam>
<lparam>Address:2997 10647</lparam>
<lparam>Address:2998 10648</lparam>
<lparam>Address:2999 10649</lparam>
<lparam>Address:3000 8192</lparam>
<lparam>Address:3001 12289</lparam>
<lparam>Address:3002 12290</lparam>
<lparam>Address:3003 12291</lparam>
<lparam>Address:3004 12292</lparam>
<lparam>Address:3005 12293</lparam>
<lparam>Address:3006 12294</lparam>
<lparam>Address:3007 12295</lparam>
<lparam>Address:3008 12296</lparam>
<lparam>Address:3009 12297</lparam>
<lparam>Address:3010 12304</lparam>
<lparam>Address:3011 12305</lparam>
<lparam>Address:3012 12306</lparam>
<lparam>Address:3013 12307</lparam>
<lparam>Address:3014 12308</lparam>
<lparam>Address:3015 12309</lparam>
<lparam>Address:3016 12310</lparam>
<lparam>Address:3017 12311</lparam>
<lparam>Address:3018 12312</lparam>
<lparam>Address:3019 12313</lparam>
<lparam>Address:3020 12320</lparam>
<lparam>Address:3021 12321</lparam>
<lparam>Address:3022 12322</lparam>
<lparam>Address:3023 12323</lparam>
<lparam>Address:3024 12324</lparam>
<lparam>Address:3025 12325</lparam>
<lparam>Address:3026 12326</lparam>
<lparam>Address:3027 12327</lparam>
<lparam>Address:3028 12328</lparam>
<lparam>Address:3029 12329</lparam>
<lparam>Address:3030 12336</lparam>
<lparam>Address:3031 12337</lparam>
<lparam>Address:3032 12338</lparam>
<lparam>Address:3033 12339</lparam>
<lparam>Address:3034 12340</lparam>
<lparam>Address:3035 12341</lparam>
<lparam>Address:3036 12342</lparam>
<lparam>Address:3037 12343</lparam>
<lparam>Address:3038 12344</lparam>
<lparam>Address:3039 12345</lparam>
<lparam>Address:3040 12352</lparam>
<lparam>Address:3041 12353</lparam>
<lparam>Address:3042 12354</lparam>
<lparam>Address:3043 12355</lparam>
<lparam>Address:3044 12356</lparam>
<lparam>Address:3045 12357</lparam>
<lparam>Address:3046 12358</lparam>
<lparam>Address:3047 12359</lparam>
<lparam>Address:3048 12360</lparam>
<lparam>Address:3049 12361</lparam>
<lparam>Address:3050 12368</lparam>
<lparam>Address:3051 12369</lparam>
<lparam>Address:3052 12370</lparam>
<lparam>Address:3053 12371</lparam>
<lparam>Address:3054 12372</lparam>
<lparam>Address:3055 12373</lparam>
<lparam>Address:3056 12374</lparam>
<lparam>Address:3057 12375</lparam>
<lparam>Address:3058 12376</lparam>
<lparam>Address:3059 12377</lparam>
<lparam>Address:3060 12384</lparam>
<lparam>Address:3061 12385</lparam>
<lparam>Address:3062 12386</lparam>
<lparam>Address:3063 12387</lparam>
<lparam>Address:3064 12388</lparam>
<lparam>Address:3065 12389</lparam>
<lparam>Address:3066 12390</lparam>
<lparam>Address:3067 12391</lparam>
<lparam>Address:3068 12392</lparam>
<lparam>Address:3069 12393</lparam>
<lparam>Address:3070 12400</lparam>
<lparam>Address:3071 12401</lparam>
<lparam>Address:3072 12402</lparam>
<lparam>Address:3073 12403</lparam>
<lparam>Address:3074 12404</lparam>
<lparam>Address:3075 12405</lparam>
<lparam>Address:3076 12406</lparam>
<lparam>Address:3077 12407</lparam>
<lparam>Address:3078 12408</lparam>
<lparam>Address:3079 12409</lparam>
<lparam>Address:3080 12416</lparam>
<lparam>Address:3081 12417</lparam>
<lparam>Address:3082 12418</lparam>
<lparam>Address:3083 12419</lparam>
<lparam>Address:3084 12420</lparam>
<lparam>Address:3085 12421</lparam>
<lparam>Address:3086 12422</lparam>
<lparam>Address:3087 12423</lparam>
<lparam>Address:3088 12424</lparam>
<lparam>Address:3089 12425</lparam>
<lparam>Address:3090 12432</lparam>
<lparam>Address:3091 12433</lparam>
<lparam>Address:3092 12434</lparam>
<lparam>Address:3093 12435</lparam>
<lparam>Address:3094 12436</lparam>
<lparam>Address:3095 12437</lparam>
<lparam>Address:3096 12438</lparam>
<lparam>Address:3097 12439</lparam>
<lparam>Address:3098 12440</lparam>
<lparam>Address:3099 12441</lparam>
<lparam>Address:3100 12544</lparam>
<lparam>Address:3101 12545</lparam>
<lparam>Address:3102 12546</lparam>
<lparam>Address:3103 12547</lparam>
<lparam>Address:3104 12548</lparam>
<lparam>Address:3105 12549</lparam>
<lparam>Address:3106 12550</lparam>
<lparam>Address:3107 12551</lparam>
<lparam>Address:3108 12552</lparam>
<lparam>Address:3109 12553</lparam>
<lparam>Address:3110 12560</lparam>
<lparam>Address:3111 12561</lparam>
<lparam>Address:3112 12562</lparam>
<lparam>Address:3113 12563</lparam>
<lparam>Address:3114 12564</lparam>
<lparam>Address:3115 12565</lparam>
<lparam>Address:3116 12566</lparam>
<lparam>Address:3117 12567</lparam>
<lparam>Address:3118 12568</lparam>
<lparam>Address:3119 12569</lparam>
<lparam>Address:3120 12576</lparam>
<lparam>Address:3121 12577</lparam>
<lparam>Address:3122 12578</lparam>
<lparam>Address:3123 12579</lparam>
<lparam>Address:3124 12580</lparam>
<lparam>Address:3125 12581</lparam>
<lparam>Address:3126 12582</lparam>
<lparam>Address:3127 12583</lparam>
<lparam>Address:3128 12584</lparam>
<lparam>Address:3129 12585</lparam>
<lparam>Address:3130 12592</lparam>
<lparam>Address:3131 12593</lparam>
<lparam>Address:3132 12594</lparam>
<lparam>Address:3133 12595</lparam>
<lparam>Address:3134 12596</lparam>
<lparam>Address:3135 12597</lparam>
<lparam>Address:3136 12598</lparam>
<lparam>Address:3137 12599</lparam>
<lparam>Address:3138 12600</lparam>
<lparam>Address:3139 12601</lparam>
<lparam>Address:3140 12608</lparam>
<lparam>Address:3141 12609</lparam>
<lparam>Address:3142 12610</lparam>
<lparam>Address:3143 12611</lparam>
<lparam>Address:3144 12612</lparam>
<lparam>Address:3145 12613</lparam>
<lparam>Address:3146 12614</lparam>
<lparam>Address:3147 12615</lparam>
<lparam>Address:3148 12616</lparam>
<lparam>Address:3149 12617</lparam>
<lparam>Address:3150 12624</lparam>
<lparam>Address:3151 12625</lparam>
<lparam>Address:3152 12626</lparam>
<lparam>Address:3153 12627</lparam>
<lparam>Address:3154 12628</lparam>
<lparam>Address:3155 12629</lparam>
<lparam>Address:3156 12630</lparam>
<lparam>Address:3157 12631</lparam>
<lparam>Address:3158 12632</lparam>
<lparam>Address:3159 12633</lparam>
<lparam>Address:3160 12640</lparam>
<lparam>Address:3161 12641</lparam>
<lparam>Address:3162 12642</lparam>
<lparam>Address:3163 12643</lparam>
<lparam>Address:3164 12644</lparam>
<lparam>Address:3165 12645</lparam>
<lparam>Address:3166 12646</lparam>
<lparam>Address:3167 12647</lparam>
<lparam>Address:3168 12648</lparam>
<lparam>Address:3169 12649</lparam>
<lparam>Address:3170 12656</lparam>
<lparam>Address:3171 12657</lparam>
<lparam>Address:3172 12658</lparam>
<lparam>Address:3173 12659</lparam>
<lparam>Address:3174 12660</lparam>
<lparam>Address:3175 12661</lparam>
<lparam>Address:3176 12662</lparam>
<lparam>Address:3177 12663</lparam>
<lparam>Address:3178 12664</lparam>
<lparam>Address:3179 12665</lparam>
<lparam>Address:3180 12672</lparam>
<lparam>Address:3181 12673</lparam>
<lparam>Address:3182 12674</lparam>
<lparam>Address:3183 12675</lparam>
<lparam>Address:3184 12676</lparam>
<lparam>Address:3185 12677</lparam>
<lparam>Address:3186 12678</lparam>
<lparam>Address:3187 12679</lparam>
<lparam>Address:3188 12680</lparam>
<lparam>Address:3189 12681</lparam>
<lparam>Address:3190 12688</lparam>
<lparam>Address:3191 12689</lparam>
<lparam>Address:3192 12690</lparam>
<lparam>Address:3193 12691</lparam>
<lparam>Address:3194 12692</lparam>
<lparam>Address:3195 12693</lparam>
<lparam>Address:3196 12694</lparam>
<lparam>Address:3197 12695</lparam>
<lparam>Address:3198 12696</lparam>
<lparam>Address:3199 12697</lparam>
<lparam>Address:3200 12800</lparam>
<lparam>Address:3201 12801</lparam>
<lparam>Address:3202 12802</lparam>
<lparam>Address:3203 12803</lparam>
<lparam>Address:3204 12804</lparam>
<lparam>Address:3205 12805</lparam>
<lparam>Address:3206 12806</lparam>
<lparam>Address:3207 12807</lparam>
<lparam>Address:3208 12808</lparam>
<lparam>Address:3209 12809</lparam>
<lparam>Address:3210 12816</lparam>
<lparam>Address:3211 12817</lparam>
<lparam>Address:3212 12818</lparam>
<lparam>Address:3213 12819</lparam>
<lparam>Address:3214 12820</lparam>
<lparam>Address:3215 12821</lparam>
<lparam>Address:3216 12822</lparam>
<lparam>Address:3217 12823</lparam>
<lparam>Address:3218 12824</lparam>
<lparam>Address:3219 12825</lparam>
<lparam>Address:3220 12832</lparam>
<lparam>Address:3221 12833</lparam>
<lparam>Address:3222 12834</lparam>
<lparam>Address:3223 12835</lparam>
<lparam>Address:3224 12836</lparam>
<lparam>Address:3225 12837</lparam>
<lparam>Address:3226 12838</lparam>
<lparam>Address:3227 12839</lparam>
<lparam>Address:3228 12840</lparam>
<lparam>Address:3229 12841</lparam>
<lparam>Address:3230 12848</lparam>
<lparam>Address:3231 12849</lparam>
<lparam>Address:3232 12850</lparam>
<lparam>Address:3233 12851</lparam>
<lparam>Address:3234 12852</lparam>
<lparam>Address:3235 12853</lparam>
<lparam>Address:3236 12854</lparam>
<lparam>Address:3237 12855</lparam>
<lparam>Address:3238 12856</lparam>
<lparam>Address:3239 12857</lparam>
<lparam>Address:3240 12864</lparam>
<lparam>Address:3241 12865</lparam>
<lparam>Address:3242 12866</lparam>
<lparam>Address:3243 12867</lparam>
<lparam>Address:3244 12868</lparam>
<lparam>Address:3245 12869</lparam>
<lparam>Address:3246 12870</lparam>
<lparam>Address:3247 12871</lparam>
<lparam>Address:3248 12872</lparam>
<lparam>Address:3249 12873</lparam>
<lparam>Address:3250 12880</lparam>
<lparam>Address:3251 12881</lparam>
<lparam>Address:3252 12882</lparam>
<lparam>Address:3253 12883</lparam>
<lparam>Address:3254 12884</lparam>
<lparam>Address:3255 12885</lparam>
<lparam>Address:3256 12886</lparam>
<lparam>Address:3257 12887</lparam>
<lparam>Address:3258 12888</lparam>
<lparam>Address:3259 12889</lparam>
<lparam>Address:3260 12896</lparam>
<lparam>Address:3261 12897</lparam>
<lparam>Address:3262 12898</lparam>
<lparam>Address:3263 12899</lparam>
<lparam>Address:3264 12900</lparam>
<lparam>Address:3265 12901</lparam>
<lparam>Address:3266 12902</lparam>
<lparam>Address:3267 12903</lparam>
<lparam>Address:3268 12904</lparam>
<lparam>Address:3269 12905</lparam>
<lparam>Address:3270 12912</lparam>
<lparam>Address:3271 12913</lparam>
<lparam>Address:3272 12914</lparam>
<lparam>Address:3273 12915</lparam>
<lparam>Address:3274 12916</lparam>
<lparam>Address:3275 12917</lparam>
<lparam>Address:3276 12918</lparam>
<lparam>Address:3277 12919</lparam>
<lparam>Address:3278 12920</lparam>
<lparam>Address:3279 12921</lparam>
<lparam>Address:3280 12928</lparam>
<lparam>Address:3281 12929</lparam>
<lparam>Address:3282 12930</lparam>
<lparam>Address:3283 12931</lparam>
<lparam>Address:3284 12932</lparam>
<lparam>Address:3285 12933</lparam>
<lparam>Address:3286 12934</lparam>
<lparam>Address:3287 12935</lparam>
<lparam>Address:3288 12936</lparam>
<lparam>Address:3289 12937</lparam>
<lparam>Address:3290 12944</lparam>
<lparam>Address:3291 12945</lparam>
<lparam>Address:3292 12946</lparam>
<lparam>Address:3293 12947</lparam>
<lparam>Address:3294 12948</lparam>
<lparam>Address:3295 12949</lparam>
<lparam>Address:3296 12950</lparam>
<lparam>Address:3297 12951</lparam>
<lparam>Address:3298 12952</lparam>
<lparam>Address:3299 12953</lparam>
<lparam>Address:3300 13056</lparam>
<lparam>Address:3301 13057</lparam>
<lparam>Address:3302 13058</lparam>
<lparam>Address:3303 13059</lparam>
<lparam>Address:3304 13060</lparam>
<lparam>Address:3305 13061</lparam>
<lparam>Address:3306 13062</lparam>
<lparam>Address:3307 13063</lparam>
<lparam>Address:3308 13064</lparam>
<lparam>Address:3309 13065</lparam>
<lparam>Address:3310 13072</lparam>
<lparam>Address:3311 13073</lparam>
<lparam>Address:3312 13074</lparam>
<lparam>Address:3313 13075</lparam>
<lparam>Address:3314 13076</lparam>
<lparam>Address:3315 13077</lparam>
<lparam>Address:3316 13078</lparam>
<lparam>Address:3317 13079</lparam>
<lparam>Address:3318 13080</lparam>
<lparam>Address:3319 13081</lparam>
<lparam>Address:3320 13088</lparam>
<lparam>Address:3321 13089</lparam>
<lparam>Address:3322 13090</lparam>
<lparam>Address:3323 13091</lparam>
<lparam>Address:3324 13092</lparam>
<lparam>Address:3325 13093</lparam>
<lparam>Address:3326 13094</lparam>
<lparam>Address:3327 13095</lparam>
<lparam>Address:3328 13096</lparam>
<lparam>Address:3329 13097</lparam>
<lparam>Address:3330 13104</lparam>
<lparam>Address:3331 13105</lparam>
<lparam>Address:3332 13106</lparam>
<lparam>Address:3333 13107</lparam>
<lparam>Address:3334 13108</lparam>
<lparam>Address:3335 13109</lparam>
<lparam>Address:3336 13110</lparam>
<lparam>Address:3337 13111</lparam>
<lparam>Address:3338 13112</lparam>
<lparam>Address:3339 13113</lparam>
<lparam>Address:3340 13120</lparam>
<lparam>Address:3341 13121</lparam>
<lparam>Address:3342 13122</lparam>
<lparam>Address:3343 13123</lparam>
<lparam>Address:3344 13124</lparam>
<lparam>Address:3345 13125</lparam>
<lparam>Address:3346 13126</lparam>
<lparam>Address:3347 13127</lparam>
<lparam>Address:3348 13128</lparam>
<lparam>Address:3349 13129</lparam>
<lparam>Address:3350 13136</lparam>
<lparam>Address:3351 13137</lparam>
<lparam>Address:3352 13138</lparam>
<lparam>Address:3353 13139</lparam>
<lparam>Address:3354 13140</lparam>
<lparam>Address:3355 13141</lparam>
<lparam>Address:3356 13142</lparam>
<lparam>Address:3357 13143</lparam>
<lparam>Address:3358 13144</lparam>
<lparam>Address:3359 13145</lparam>
<lparam>Address:3360 13152</lparam>
<lparam>Address:3361 13153</lparam>
<lparam>Address:3362 13154</lparam>
<lparam>Address:3363 13155</lparam>
<lparam>Address:3364 13156</lparam>
<lparam>Address:3365 13157</lparam>
<lparam>Address:3366 13158</lparam>
<lparam>Address:3367 13159</lparam>
<lparam>Address:3368 13160</lparam>
<lparam>Address:3369 13161</lparam>
<lparam>Address:3370 13168</lparam>
<lparam>Address:3371 13169</lparam>
<lparam>Address:3372 13170</lparam>
<lparam>Address:3373 13171</lparam>
<lparam>Address:3374 13172</lparam>
<lparam>Address:3375 13173</lparam>
<lparam>Address:3376 13174</lparam>
<lparam>Address:3377 13175</lparam>
<lparam>Address:3378 13176</lparam>
<lparam>Address:3379 13177</lparam>
<lparam>Address:3380 13184</lparam>
<lparam>Address:3381 13185</lparam>
<lparam>Address:3382 13186</lparam>
<lparam>Address:3383 13187</lparam>
<lparam>Address:3384 13188</lparam>
<lparam>Address:3385 13189</lparam>
<lparam>Address:3386 13190</lparam>
<lparam>Address:3387 13191</lparam>
<lparam>Address:3388 13192</lparam>
<lparam>Address:3389 13193</lparam>
<lparam>Address:3390 13200</lparam>
<lparam>Address:3391 13201</lparam>
<lparam>Address:3392 13202</lparam>
<lparam>Address:3393 13203</lparam>
<lparam>Address:3394 13204</lparam>
<lparam>Address:3395 13205</lparam>
<lparam>Address:3396 13206</lparam>
<lparam>Address:3397 13207</lparam>
<lparam>Address:3398 13208</lparam>
<lparam>Address:3399 13209</lparam>
<lparam>Address:3400 13312</lparam>
<lparam>Address:3401 13313</lparam>
<lparam>Address:3402 13314</lparam>
<lparam>Address:3403 13315</lparam>
<lparam>Address:3404 13316</lparam>
<lparam>Address:3405 13317</lparam>
<lparam>Address:3406 13318</lparam>
<lparam>Address:3407 13319</lparam>
<lparam>Address:3408 13320</lparam>
<lparam>Address:3409 13321</lparam>
<lparam>Address:3410 13328</lparam>
<lparam>Address:3411 13329</lparam>
<lparam>Address:3412 13330</lparam>
<lparam>Address:3413 13331</lparam>
<lparam>Address:3414 13332</lparam>
<lparam>Address:3415 13333</lparam>
<lparam>Address:3416 13334</lparam>
<lparam>Address:3417 13335</lparam>
<lparam>Address:3418 13336</lparam>
<lparam>Address:3419 13337</lparam>
<lparam>Address:3420 13344</lparam>
<lparam>Address:3421 13345</lparam>
<lparam>Address:3422 13346</lparam>
<lparam>Address:3423 13347</lparam>
<lparam>Address:3424 13348</lparam>
<lparam>Address:3425 13349</lparam>
<lparam>Address:3426 13350</lparam>
<lparam>Address:3427 13351</lparam>
<lparam>Address:3428 13352</lparam>
<lparam>Address:3429 13353</lparam>
<lparam>Address:3430 13360</lparam>
<lparam>Address:3431 13361</lparam>
<lparam>Address:3432 13362</lparam>
<lparam>Address:3433 13363</lparam>
<lparam>Address:3434 13364</lparam>
<lparam>Address:3435 13365</lparam>
<lparam>Address:3436 13366</lparam>
<lparam>Address:3437 13367</lparam>
<lparam>Address:3438 13368</lparam>
<lparam>Address:3439 13369</lparam>
<lparam>Address:3440 13376</lparam>
<lparam>Address:3441 13377</lparam>
<lparam>Address:3442 13378</lparam>
<lparam>Address:3443 13379</lparam>
<lparam>Address:3444 13380</lparam>
<lparam>Address:3445 13381</lparam>
<lparam>Address:3446 13382</lparam>
<lparam>Address:3447 13383</lparam>
<lparam>Address:3448 13384</lparam>
<lparam>Address:3449 13385</lparam>
<lparam>Address:3450 13392</lparam>
<lparam>Address:3451 13393</lparam>
<lparam>Address:3452 13394</lparam>
<lparam>Address:3453 13395</lparam>
<lparam>Address:3454 13396</lparam>
<lparam>Address:3455 13397</lparam>
<lparam>Address:3456 13398</lparam>
<lparam>Address:3457 13399</lparam>
<lparam>Address:3458 13400</lparam>
<lparam>Address:3459 13401</lparam>
<lparam>Address:3460 13408</lparam>
<lparam>Address:3461 13409</lparam>
<lparam>Address:3462 13410</lparam>
<lparam>Address:3463 13411</lparam>
<lparam>Address:3464 13412</lparam>
<lparam>Address:3465 13413</lparam>
<lparam>Address:3466 13414</lparam>
<lparam>Address:3467 13415</lparam>
<lparam>Address:3468 13416</lparam>
<lparam>Address:3469 13417</lparam>
<lparam>Address:3470 13424</lparam>
<lparam>Address:3471 13425</lparam>
<lparam>Address:3472 13426</lparam>
<lparam>Address:3473 13427</lparam>
<lparam>Address:3474 13428</lparam>
<lparam>Address:3475 13429</lparam>
<lparam>Address:3476 13430</lparam>
<lparam>Address:3477 13431</lparam>
<lparam>Address:3478 13432</lparam>
<lparam>Address:3479 13433</lparam>
<lparam>Address:3480 13440</lparam>
<lparam>Address:3481 13441</lparam>
<lparam>Address:3482 13442</lparam>
<lparam>Address:3483 13443</lparam>
<lparam>Address:3484 13444</lparam>
<lparam>Address:3485 13445</lparam>
<lparam>Address:3486 13446</lparam>
<lparam>Address:3487 13447</lparam>
<lparam>Address:3488 13448</lparam>
<lparam>Address:3489 13449</lparam>
<lparam>Address:3490 13456</lparam>
<lparam>Address:3491 13457</lparam>
<lparam>Address:3492 13458</lparam>
<lparam>Address:3493 13459</lparam>
<lparam>Address:3494 13460</lparam>
<lparam>Address:3495 13461</lparam>
<lparam>Address:3496 13462</lparam>
<lparam>Address:3497 13463</lparam>
<lparam>Address:3498 13464</lparam>
<lparam>Address:3499 13465</lparam>
<lparam>Address:3500 13568</lparam>
<lparam>Address:3501 13569</lparam>
<lparam>Address:3502 13570</lparam>
<lparam>Address:3503 13571</lparam>
<lparam>Address:3504 13572</lparam>
<lparam>Address:3505 13573</lparam>
<lparam>Address:3506 13574</lparam>
<lparam>Address:3507 13575</lparam>
<lparam>Address:3508 13576</lparam>
<lparam>Address:3509 13577</lparam>
<lparam>Address:3510 13584</lparam>
<lparam>Address:3511 13585</lparam>
<lparam>Address:3512 13586</lparam>
<lparam>Address:3513 13587</lparam>
<lparam>Address:3514 13588</lparam>
<lparam>Address:3515 13589</lparam>
<lparam>Address:3516 13590</lparam>
<lparam>Address:3517 13591</lparam>
<lparam>Address:3518 13592</lparam>
<lparam>Address:3519 13593</lparam>
<lparam>Address:3520 13600</lparam>
<lparam>Address:3521 13601</lparam>
<lparam>Address:3522 13602</lparam>
<lparam>Address:3523 13603</lparam>
<lparam>Address:3524 13604</lparam>
<lparam>Address:3525 13605</lparam>
<lparam>Address:3526 13606</lparam>
<lparam>Address:3527 13607</lparam>
<lparam>Address:3528 13608</lparam>
<lparam>Address:3529 13609</lparam>
<lparam>Address:3530 13616</lparam>
<lparam>Address:3531 13617</lparam>
<lparam>Address:3532 13618</lparam>
<lparam>Address:3533 13619</lparam>
<lparam>Address:3534 13620</lparam>
<lparam>Address:3535 13621</lparam>
<lparam>Address:3536 13622</lparam>
<lparam>Address:3537 13623</lparam>
<lparam>Address:3538 13624</lparam>
<lparam>Address:3539 13625</lparam>
<lparam>Address:3540 13632</lparam>
<lparam>Address:3541 13633</lparam>
<lparam>Address:3542 13634</lparam>
<lparam>Address:3543 13635</lparam>
<lparam>Address:3544 13636</lparam>
<lparam>Address:3545 13637</lparam>
<lparam>Address:3546 13638</lparam>
<lparam>Address:3547 13639</lparam>
<lparam>Address:3548 13640</lparam>
<lparam>Address:3549 13641</lparam>
<lparam>Address:3550 13648</lparam>
<lparam>Address:3551 13649</lparam>
<lparam>Address:3552 13650</lparam>
<lparam>Address:3553 13651</lparam>
<lparam>Address:3554 13652</lparam>
<lparam>Address:3555 13653</lparam>
<lparam>Address:3556 13654</lparam>
<lparam>Address:3557 13655</lparam>
<lparam>Address:3558 13656</lparam>
<lparam>Address:3559 13657</lparam>
<lparam>Address:3560 13664</lparam>
<lparam>Address:3561 13665</lparam>
<lparam>Address:3562 13666</lparam>
<lparam>Address:3563 13667</lparam>
<lparam>Address:3564 13668</lparam>
<lparam>Address:3565 13669</lparam>
<lparam>Address:3566 13670</lparam>
<lparam>Address:3567 13671</lparam>
<lparam>Address:3568 13672</lparam>
<lparam>Address:3569 13673</lparam>
<lparam>Address:3570 13680</lparam>
<lparam>Address:3571 13681</lparam>
<lparam>Address:3572 13682</lparam>
<lparam>Address:3573 13683</lparam>
<lparam>Address:3574 13684</lparam>
<lparam>Address:3575 13685</lparam>
<lparam>Address:3576 13686</lparam>
<lparam>Address:3577 13687</lparam>
<lparam>Address:3578 13688</lparam>
<lparam>Address:3579 13689</lparam>
<lparam>Address:3580 13696</lparam>
<lparam>Address:3581 13697</lparam>
<lparam>Address:3582 13698</lparam>
<lparam>Address:3583 13699</lparam>
<lparam>Address:3584 13700</lparam>
<lparam>Address:3585 13701</lparam>
<lparam>Address:3586 13702</lparam>
<lparam>Address:3587 13703</lparam>
<lparam>Address:3588 13704</lparam>
<lparam>Address:3589 13705</lparam>
<lparam>Address:3590 13712</lparam>
<lparam>Address:3591 13713</lparam>
<lparam>Address:3592 13714</lparam>
<lparam>Address:3593 13715</lparam>
<lparam>Address:3594 13716</lparam>
<lparam>Address:3595 13717</lparam>
<lparam>Address:3596 13718</lparam>
<lparam>Address:3597 13719</lparam>
<lparam>Address:3598 13720</lparam>
<lparam>Address:3599 13721</lparam>
<lparam>Address:3600 13824</lparam>
<lparam>Address:3601 13825</lparam>
<lparam>Address:3602 13826</lparam>
<lparam>Address:3603 13827</lparam>
<lparam>Address:3604 13828</lparam>
<lparam>Address:3605 13829</lparam>
<lparam>Address:3606 13830</lparam>
<lparam>Address:3607 13831</lparam>
<lparam>Address:3608 13832</lparam>
<lparam>Address:3609 13833</lparam>
<lparam>Address:3610 13840</lparam>
<lparam>Address:3611 13841</lparam>
<lparam>Address:3612 13842</lparam>
<lparam>Address:3613 13843</lparam>
<lparam>Address:3614 13844</lparam>
<lparam>Address:3615 13845</lparam>
<lparam>Address:3616 13846</lparam>
<lparam>Address:3617 13847</lparam>
<lparam>Address:3618 13848</lparam>
<lparam>Address:3619 13849</lparam>
<lparam>Address:3620 13856</lparam>
<lparam>Address:3621 13857</lparam>
<lparam>Address:3622 13858</lparam>
<lparam>Address:3623 13859</lparam>
<lparam>Address:3624 13860</lparam>
<lparam>Address:3625 13861</lparam>
<lparam>Address:3626 13862</lparam>
<lparam>Address:3627 13863</lparam>
<lparam>Address:3628 13864</lparam>
<lparam>Address:3629 13865</lparam>
<lparam>Address:3630 13872</lparam>
<lparam>Address:3631 13873</lparam>
<lparam>Address:3632 13874</lparam>
<lparam>Address:3633 13875</lparam>
<lparam>Address:3634 13876</lparam>
<lparam>Address:3635 13877</lparam>
<lparam>Address:3636 13878</lparam>
<lparam>Address:3637 13879</lparam>
<lparam>Address:3638 13880</lparam>
<lparam>Address:3639 13881</lparam>
<lparam>Address:3640 13888</lparam>
<lparam>Address:3641 13889</lparam>
<lparam>Address:3642 13890</lparam>
<lparam>Address:3643 13891</lparam>
<lparam>Address:3644 13892</lparam>
<lparam>Address:3645 13893</lparam>
<lparam>Address:3646 13894</lparam>
<lparam>Address:3647 13895</lparam>
<lparam>Address:3648 13896</lparam>
<lparam>Address:3649 13897</lparam>
<lparam>Address:3650 13904</lparam>
<lparam>Address:3651 13905</lparam>
<lparam>Address:3652 13906</lparam>
<lparam>Address:3653 13907</lparam>
<lparam>Address:3654 13908</lparam>
<lparam>Address:3655 13909</lparam>
<lparam>Address:3656 13910</lparam>
<lparam>Address:3657 13911</lparam>
<lparam>Address:3658 13912</lparam>
<lparam>Address:3659 13913</lparam>
<lparam>Address:3660 13920</lparam>
<lparam>Address:3661 13921</lparam>
<lparam>Address:3662 13922</lparam>
<lparam>Address:3663 13923</lparam>
<lparam>Address:3664 13924</lparam>
<lparam>Address:3665 13925</lparam>
<lparam>Address:3666 13926</lparam>
<lparam>Address:3667 13927</lparam>
<lparam>Address:3668 13928</lparam>
<lparam>Address:3669 13929</lparam>
<lparam>Address:3670 13936</lparam>
<lparam>Address:3671 13937</lparam>
<lparam>Address:3672 13938</lparam>
<lparam>Address:3673 13939</lparam>
<lparam>Address:3674 13940</lparam>
<lparam>Address:3675 13941</lparam>
<lparam>Address:3676 13942</lparam>
<lparam>Address:3677 13943</lparam>
<lparam>Address:3678 13944</lparam>
<lparam>Address:3679 13945</lparam>
<lparam>Address:3680 13952</lparam>
<lparam>Address:3681 13953</lparam>
<lparam>Address:3682 13954</lparam>
<lparam>Address:3683 13955</lparam>
<lparam>Address:3684 13956</lparam>
<lparam>Address:3685 13957</lparam>
<lparam>Address:3686 13958</lparam>
<lparam>Address:3687 13959</lparam>
<lparam>Address:3688 13960</lparam>
<lparam>Address:3689 13961</lparam>
<lparam>Address:3690 13968</lparam>
<lparam>Address:3691 13969</lparam>
<lparam>Address:3692 13970</lparam>
<lparam>Address:3693 13971</lparam>
<lparam>Address:3694 13972</lparam>
<lparam>Address:3695 13973</lparam>
<lparam>Address:3696 13974</lparam>
<lparam>Address:3697 13975</lparam>
<lparam>Address:3698 13976</lparam>
<lparam>Address:3699 13977</lparam>
<lparam>Address:3700 14080</lparam>
<lparam>Address:3701 14081</lparam>
<lparam>Address:3702 14082</lparam>
<lparam>Address:3703 14083</lparam>
<lparam>Address:3704 14084</lparam>
<lparam>Address:3705 14085</lparam>
<lparam>Address:3706 14086</lparam>
<lparam>Address:3707 14087</lparam>
<lparam>Address:3708 14088</lparam>
<lparam>Address:3709 14089</lparam>
<lparam>Address:3710 14096</lparam>
<lparam>Address:3711 14097</lparam>
<lparam>Address:3712 14098</lparam>
<lparam>Address:3713 14099</lparam>
<lparam>Address:3714 14100</lparam>
<lparam>Address:3715 14101</lparam>
<lparam>Address:3716 14102</lparam>
<lparam>Address:3717 14103</lparam>
<lparam>Address:3718 14104</lparam>
<lparam>Address:3719 14105</lparam>
<lparam>Address:3720 14112</lparam>
<lparam>Address:3721 14113</lparam>
<lparam>Address:3722 14114</lparam>
<lparam>Address:3723 14115</lparam>
<lparam>Address:3724 14116</lparam>
<lparam>Address:3725 14117</lparam>
<lparam>Address:3726 14118</lparam>
<lparam>Address:3727 14119</lparam>
<lparam>Address:3728 14120</lparam>
<lparam>Address:3729 14121</lparam>
<lparam>Address:3730 14128</lparam>
<lparam>Address:3731 14129</lparam>
<lparam>Address:3732 14130</lparam>
<lparam>Address:3733 14131</lparam>
<lparam>Address:3734 14132</lparam>
<lparam>Address:3735 14133</lparam>
<lparam>Address:3736 14134</lparam>
<lparam>Address:3737 14135</lparam>
<lparam>Address:3738 14136</lparam>
<lparam>Address:3739 14137</lparam>
<lparam>Address:3740 14144</lparam>
<lparam>Address:3741 14145</lparam>
<lparam>Address:3742 14146</lparam>
<lparam>Address:3743 14147</lparam>
<lparam>Address:3744 14148</lparam>
<lparam>Address:3745 14149</lparam>
<lparam>Address:3746 14150</lparam>
<lparam>Address:3747 14151</lparam>
<lparam>Address:3748 14152</lparam>
<lparam>Address:3749 14153</lparam>
<lparam>Address:3750 14160</lparam>
<lparam>Address:3751 14161</lparam>
<lparam>Address:3752 14162</lparam>
<lparam>Address:3753 14163</lparam>
<lparam>Address:3754 14164</lparam>
<lparam>Address:3755 14165</lparam>
<lparam>Address:3756 14166</lparam>
<lparam>Address:3757 14167</lparam>
<lparam>Address:3758 14168</lparam>
<lparam>Address:3759 14169</lparam>
<lparam>Address:3760 14176</lparam>
<lparam>Address:3761 14177</lparam>
<lparam>Address:3762 14178</lparam>
<lparam>Address:3763 14179</lparam>
<lparam>Address:3764 14180</lparam>
<lparam>Address:3765 14181</lparam>
<lparam>Address:3766 14182</lparam>
<lparam>Address:3767 14183</lparam>
<lparam>Address:3768 14184</lparam>
<lparam>Address:3769 14185</lparam>
<lparam>Address:3770 14192</lparam>
<lparam>Address:3771 14193</lparam>
<lparam>Address:3772 14194</lparam>
<lparam>Address:3773 14195</lparam>
<lparam>Address:3774 14196</lparam>
<lparam>Address:3775 14197</lparam>
<lparam>Address:3776 14198</lparam>
<lparam>Address:3777 14199</lparam>
<lparam>Address:3778 14200</lparam>
<lparam>Address:3779 14201</lparam>
<lparam>Address:3780 14208</lparam>
<lparam>Address:3781 14209</lparam>
<lparam>Address:3782 14210</lparam>
<lparam>Address:3783 14211</lparam>
<lparam>Address:3784 14212</lparam>
<lparam>Address:3785 14213</lparam>
<lparam>Address:3786 14214</lparam>
<lparam>Address:3787 14215</lparam>
<lparam>Address:3788 14216</lparam>
<lparam>Address:3789 14217</lparam>
<lparam>Address:3790 14224</lparam>
<lparam>Address:3791 14225</lparam>
<lparam>Address:3792 14226</lparam>
<lparam>Address:3793 14227</lparam>
<lparam>Address:3794 14228</lparam>
<lparam>Address:3795 14229</lparam>
<lparam>Address:3796 14230</lparam>
<lparam>Address:3797 14231</lparam>
<lparam>Address:3798 14232</lparam>
<lparam>Address:3799 14233</lparam>
<lparam>Address:3800 14336</lparam>
<lparam>Address:3801 14337</lparam>
<lparam>Address:3802 14338</lparam>
<lparam>Address:3803 14339</lparam>
<lparam>Address:3804 14340</lparam>
<lparam>Address:3805 14341</lparam>
<lparam>Address:3806 14342</lparam>
<lparam>Address:3807 14343</lparam>
<lparam>Address:3808 14344</lparam>
<lparam>Address:3809 14345</lparam>
<lparam>Address:3810 14352</lparam>
<lparam>Address:3811 14353</lparam>
<lparam>Address:3812 14354</lparam>
<lparam>Address:3813 14355</lparam>
<lparam>Address:3814 14356</lparam>
<lparam>Address:3815 14357</lparam>
<lparam>Address:3816 14358</lparam>
<lparam>Address:3817 14359</lparam>
<lparam>Address:3818 14360</lparam>
<lparam>Address:3819 14361</lparam>
<lparam>Address:3820 14368</lparam>
<lparam>Address:3821 14369</lparam>
<lparam>Address:3822 14370</lparam>
<lparam>Address:3823 14371</lparam>
<lparam>Address:3824 14372</lparam>
<lparam>Address:3825 14373</lparam>
<lparam>Address:3826 14374</lparam>
<lparam>Address:3827 14375</lparam>
<lparam>Address:3828 14376</lparam>
<lparam>Address:3829 14377</lparam>
<lparam>Address:3830 14384</lparam>
<lparam>Address:3831 14385</lparam>
<lparam>Address:3832 14386</lparam>
<lparam>Address:3833 14387</lparam>
<lparam>Address:3834 14388</lparam>
<lparam>Address:3835 14389</lparam>
<lparam>Address:3836 14390</lparam>
<lparam>Address:3837 14391</lparam>
<lparam>Address:3838 14392</lparam>
<lparam>Address:3839 14393</lparam>
<lparam>Address:3840 14400</lparam>
<lparam>Address:3841 14401</lparam>
<lparam>Address:3842 14402</lparam>
<lparam>Address:3843 14403</lparam>
<lparam>Address:3844 14404</lparam>
<lparam>Address:3845 14405</lparam>
<lparam>Address:3846 14406</lparam>
<lparam>Address:3847 14407</lparam>
<lparam>Address:3848 14408</lparam>
<lparam>Address:3849 14409</lparam>
<lparam>Address:3850 14416</lparam>
<lparam>Address:3851 14417</lparam>
<lparam>Address:3852 14418</lparam>
<lparam>Address:3853 14419</lparam>
<lparam>Address:3854 14420</lparam>
<lparam>Address:3855 14421</lparam>
<lparam>Address:3856 14422</lparam>
<lparam>Address:3857 14423</lparam>
<lparam>Address:3858 14424</lparam>
<lparam>Address:3859 14425</lparam>
<lparam>Address:3860 14432</lparam>
<lparam>Address:3861 14433</lparam>
<lparam>Address:3862 14434</lparam>
<lparam>Address:3863 14435</lparam>
<lparam>Address:3864 14436</lparam>
<lparam>Address:3865 14437</lparam>
<lparam>Address:3866 14438</lparam>
<lparam>Address:3867 14439</lparam>
<lparam>Address:3868 14440</lparam>
<lparam>Address:3869 14441</lparam>
<lparam>Address:3870 14448</lparam>
<lparam>Address:3871 14449</lparam>
<lparam>Address:3872 14450</lparam>
<lparam>Address:3873 14451</lparam>
<lparam>Address:3874 14452</lparam>
<lparam>Address:3875 14453</lparam>
<lparam>Address:3876 14454</lparam>
<lparam>Address:3877 14455</lparam>
<lparam>Address:3878 14456</lparam>
<lparam>Address:3879 14457</lparam>
<lparam>Address:3880 14464</lparam>
<lparam>Address:3881 14465</lparam>
<lparam>Address:3882 14466</lparam>
<lparam>Address:3883 14467</lparam>
<lparam>Address:3884 14468</lparam>
<lparam>Address:3885 14469</lparam>
<lparam>Address:3886 14470</lparam>
<lparam>Address:3887 14471</lparam>
<lparam>Address:3888 14472</lparam>
<lparam>Address:3889 14473</lparam>
<lparam>Address:3890 14480</lparam>
<lparam>Address:3891 14481</lparam>
<lparam>Address:3892 14482</lparam>
<lparam>Address:3893 14483</lparam>
<lparam>Address:3894 14484</lparam>
<lparam>Address:3895 14485</lparam>
<lparam>Address:3896 14486</lparam>
<lparam>Address:3897 14487</lparam>
<lparam>Address:3898 14488</lparam>
<lparam>Address:3899 14489</lparam>
<lparam>Address:3900 14592</lparam>
<lparam>Address:3901 14593</lparam>
<lparam>Address:3902 14594</lparam>
<lparam>Address:3903 14595</lparam>
<lparam>Address:3904 14596</lparam>
<lparam>Address:3905 14597</lparam>
<lparam>Address:3906 14598</lparam>
<lparam>Address:3907 14599</lparam>
<lparam>Address:3908 14600</lparam>
<lparam>Address:3909 14601</lparam>
<lparam>Address:3910 14608</lparam>
<lparam>Address:3911 14609</lparam>
<lparam>Address:3912 14610</lparam>
<lparam>Address:3913 14611</lparam>
<lparam>Address:3914 14612</lparam>
<lparam>Address:3915 14613</lparam>
<lparam>Address:3916 14614</lparam>
<lparam>Address:3917 14615</lparam>
<lparam>Address:3918 14616</lparam>
<lparam>Address:3919 14617</lparam>
<lparam>Address:3920 14624</lparam>
<lparam>Address:3921 14625</lparam>
<lparam>Address:3922 14626</lparam>
<lparam>Address:3923 14627</lparam>
<lparam>Address:3924 14628</lparam>
<lparam>Address:3925 14629</lparam>
<lparam>Address:3926 14630</lparam>
<lparam>Address:3927 14631</lparam>
<lparam>Address:3928 14632</lparam>
<lparam>Address:3929 14633</lparam>
<lparam>Address:3930 14640</lparam>
<lparam>Address:3931 14641</lparam>
<lparam>Address:3932 14642</lparam>
<lparam>Address:3933 14643</lparam>
<lparam>Address:3934 14644</lparam>
<lparam>Address:3935 14645</lparam>
<lparam>Address:3936 14646</lparam>
<lparam>Address:3937 14647</lparam>
<lparam>Address:3938 14648</lparam>
<lparam>Address:3939 14649</lparam>
<lparam>Address:3940 14656</lparam>
<lparam>Address:3941 14657</lparam>
<lparam>Address:3942 14658</lparam>
<lparam>Address:3943 14659</lparam>
<lparam>Address:3944 14660</lparam>
<lparam>Address:3945 14661</lparam>
<lparam>Address:3946 14662</lparam>
<lparam>Address:3947 14663</lparam>
<lparam>Address:3948 14664</lparam>
<lparam>Address:3949 14665</lparam>
<lparam>Address:3950 14672</lparam>
<lparam>Address:3951 14673</lparam>
<lparam>Address:3952 14674</lparam>
<lparam>Address:3953 14675</lparam>
<lparam>Address:3954 14676</lparam>
<lparam>Address:3955 14677</lparam>
<lparam>Address:3956 14678</lparam>
<lparam>Address:3957 14679</lparam>
<lparam>Address:3958 14680</lparam>
<lparam>Address:3959 14681</lparam>
<lparam>Address:3960 14688</lparam>
<lparam>Address:3961 14689</lparam>
<lparam>Address:3962 14690</lparam>
<lparam>Address:3963 14691</lparam>
<lparam>Address:3964 14692</lparam>
<lparam>Address:3965 14693</lparam>
<lparam>Address:3966 14694</lparam>
<lparam>Address:3967 14695</lparam>
<lparam>Address:3968 14696</lparam>
<lparam>Address:3969 14697</lparam>
<lparam>Address:3970 14704</lparam>
<lparam>Address:3971 14705</lparam>
<lparam>Address:3972 14706</lparam>
<lparam>Address:3973 14707</lparam>
<lparam>Address:3974 14708</lparam>
<lparam>Address:3975 14709</lparam>
<lparam>Address:3976 14710</lparam>
<lparam>Address:3977 14711</lparam>
<lparam>Address:3978 14712</lparam>
<lparam>Address:3979 14713</lparam>
<lparam>Address:3980 14720</lparam>
<lparam>Address:3981 14721</lparam>
<lparam>Address:3982 14722</lparam>
<lparam>Address:3983 14723</lparam>
<lparam>Address:3984 14724</lparam>
<lparam>Address:3985 14725</lparam>
<lparam>Address:3986 14726</lparam>
<lparam>Address:3987 14727</lparam>
<lparam>Address:3988 14728</lparam>
<lparam>Address:3989 14729</lparam>
<lparam>Address:3990 14736</lparam>
<lparam>Address:3991 14737</lparam>
<lparam>Address:3992 14738</lparam>
<lparam>Address:3993 14739</lparam>
<lparam>Address:3994 14740</lparam>
<lparam>Address:3995 14741</lparam>
<lparam>Address:3996 14742</lparam>
<lparam>Address:3997 14743</lparam>
<lparam>Address:3998 14744</lparam>
<lparam>Address:3999 14745</lparam>
<lparam>Address:4000 12288</lparam>
<lparam>Address:4001 16385</lparam>
<lparam>Address:4002 16386</lparam>
<lparam>Address:4003 16387</lparam>
<lparam>Address:4004 16388</lparam>
<lparam>Address:4005 16389</lparam>
<lparam>Address:4006 16390</lparam>
<lparam>Address:4007 16391</lparam>
<lparam>Address:4008 16392</lparam>
<lparam>Address:4009 16393</lparam>
<lparam>Address:4010 16400</lparam>
<lparam>Address:4011 16401</lparam>
<lparam>Address:4012 16402</lparam>
<lparam>Address:4013 16403</lparam>
<lparam>Address:4014 16404</lparam>
<lparam>Address:4015 16405</lparam>
<lparam>Address:4016 16406</lparam>
<lparam>Address:4017 16407</lparam>
<lparam>Address:4018 16408</lparam>
<lparam>Address:4019 16409</lparam>
<lparam>Address:4020 16416</lparam>
<lparam>Address:4021 16417</lparam>
<lparam>Address:4022 16418</lparam>
<lparam>Address:4023 16419</lparam>
<lparam>Address:4024 16420</lparam>
<lparam>Address:4025 16421</lparam>
<lparam>Address:4026 16422</lparam>
<lparam>Address:4027 16423</lparam>
<lparam>Address:4028 16424</lparam>
<lparam>Address:4029 16425</lparam>
<lparam>Address:4030 16432</lparam>
<lparam>Address:4031 16433</lparam>
<lparam>Address:4032 16434</lparam>
<lparam>Address:4033 16435</lparam>
<lparam>Address:4034 16436</lparam>
<lparam>Address:4035 16437</lparam>
<lparam>Address:4036 16438</lparam>
<lparam>Address:4037 16439</lparam>
<lparam>Address:4038 16440</lparam>
<lparam>Address:4039 16441</lparam>
<lparam>Address:4040 16448</lparam>
<lparam>Address:4041 16449</lparam>
<lparam>Address:4042 16450</lparam>
<lparam>Address:4043 16451</lparam>
<lparam>Address:4044 16452</lparam>
<lparam>Address:4045 16453</lparam>
<lparam>Address:4046 16454</lparam>
<lparam>Address:4047 16455</lparam>
<lparam>Address:4048 16456</lparam>
<lparam>Address:4049 16457</lparam>
<lparam>Address:4050 16464</lparam>
<lparam>Address:4051 16465</lparam>
<lparam>Address:4052 16466</lparam>
<lparam>Address:4053 16467</lparam>
<lparam>Address:4054 16468</lparam>
<lparam>Address:4055 16469</lparam>
<lparam>Address:4056 16470</lparam>
<lparam>Address:4057 16471</lparam>
<lparam>Address:4058 16472</lparam>
<lparam>Address:4059 16473</lparam>
<lparam>Address:4060 16480</lparam>
<lparam>Address:4061 16481</lparam>
<lparam>Address:4062 16482</lparam>
<lparam>Address:4063 16483</lparam>
<lparam>Address:4064 16484</lparam>
<lparam>Address:4065 16485</lparam>
<lparam>Address:4066 16486</lparam>
<lparam>Address:4067 16487</lparam>
<lparam>Address:4068 16488</lparam>
<lparam>Address:4069 16489</lparam>
<lparam>Address:4070 16496</lparam>
<lparam>Address:4071 16497</lparam>
<lparam>Address:4072 16498</lparam>
<lparam>Address:4073 16499</lparam>
<lparam>Address:4074 16500</lparam>
<lparam>Address:4075 16501</lparam>
<lparam>Address:4076 16502</lparam>
<lparam>Address:4077 16503</lparam>
<lparam>Address:4078 16504</lparam>
<lparam>Address:4079 16505</lparam>
<lparam>Address:4080 16512</lparam>
<lparam>Address:4081 16513</lparam>
<lparam>Address:4082 16514</lparam>
<lparam>Address:4083 16515</lparam>
<lparam>Address:4084 16516</lparam>
<lparam>Address:4085 16517</lparam>
<lparam>Address:4086 16518</lparam>
<lparam>Address:4087 16519</lparam>
<lparam>Address:4088 16520</lparam>
<lparam>Address:4089 16521</lparam>
<lparam>Address:4090 16528</lparam>
<lparam>Address:4091 16529</lparam>
<lparam>Address:4092 16530</lparam>
<lparam>Address:4093 16531</lparam>
<lparam>Address:4094 16532</lparam>
<lparam>Address:4095 16533</lparam>
<lparam>Address:4096 16534</lparam>
<lparam>Address:4097 16535</lparam>
<lparam>Address:4098 16536</lparam>
<lparam>Address:4099 16537</lparam>
<lparam>Address:4100 16640</lparam>
<lparam>Address:4101 16641</lparam>
<lparam>Address:4102 16642</lparam>
<lparam>Address:4103 16643</lparam>
<lparam>Address:4104 16644</lparam>
<lparam>Address:4105 16645</lparam>
<lparam>Address:4106 16646</lparam>
<lparam>Address:4107 16647</lparam>
<lparam>Address:4108 16648</lparam>
<lparam>Address:4109 16649</lparam>
<lparam>Address:4110 16656</lparam>
<lparam>Address:4111 16657</lparam>
<lparam>Address:4112 16658</lparam>
<lparam>Address:4113 16659</lparam>
<lparam>Address:4114 16660</lparam>
<lparam>Address:4115 16661</lparam>
<lparam>Address:4116 16662</lparam>
<lparam>Address:4117 16663</lparam>
<lparam>Address:4118 16664</lparam>
<lparam>Address:4119 16665</lparam>
<lparam>Address:4120 16672</lparam>
<lparam>Address:4121 16673</lparam>
<lparam>Address:4122 16674</lparam>
<lparam>Address:4123 16675</lparam>
<lparam>Address:4124 16676</lparam>
<lparam>Address:4125 16677</lparam>
<lparam>Address:4126 16678</lparam>
<lparam>Address:4127 16679</lparam>
<lparam>Address:4128 16680</lparam>
<lparam>Address:4129 16681</lparam>
<lparam>Address:4130 16688</lparam>
<lparam>Address:4131 16689</lparam>
<lparam>Address:4132 16690</lparam>
<lparam>Address:4133 16691</lparam>
<lparam>Address:4134 16692</lparam>
<lparam>Address:4135 16693</lparam>
<lparam>Address:4136 16694</lparam>
<lparam>Address:4137 16695</lparam>
<lparam>Address:4138 16696</lparam>
<lparam>Address:4139 16697</lparam>
<lparam>Address:4140 16704</lparam>
<lparam>Address:4141 16705</lparam>
<lparam>Address:4142 16706</lparam>
<lparam>Address:4143 16707</lparam>
<lparam>Address:4144 16708</lparam>
<lparam>Address:4145 16709</lparam>
<lparam>Address:4146 16710</lparam>
<lparam>Address:4147 16711</lparam>
<lparam>Address:4148 16712</lparam>
<lparam>Address:4149 16713</lparam>
<lparam>Address:4150 16720</lparam>
<lparam>Address:4151 16721</lparam>
<lparam>Address:4152 16722</lparam>
<lparam>Address:4153 16723</lparam>
<lparam>Address:4154 16724</lparam>
<lparam>Address:4155 16725</lparam>
<lparam>Address:4156 16726</lparam>
<lparam>Address:4157 16727</lparam>
<lparam>Address:4158 16728</lparam>
<lparam>Address:4159 16729</lparam>
<lparam>Address:4160 16736</lparam>
<lparam>Address:4161 16737</lparam>
<lparam>Address:4162 16738</lparam>
<lparam>Address:4163 16739</lparam>
<lparam>Address:4164 16740</lparam>
<lparam>Address:4165 16741</lparam>
<lparam>Address:4166 16742</lparam>
<lparam>Address:4167 16743</lparam>
<lparam>Address:4168 16744</lparam>
<lparam>Address:4169 16745</lparam>
<lparam>Address:4170 16752</lparam>
<lparam>Address:4171 16753</lparam>
<lparam>Address:4172 16754</lparam>
<lparam>Address:4173 16755</lparam>
<lparam>Address:4174 16756</lparam>
<lparam>Address:4175 16757</lparam>
<lparam>Address:4176 16758</lparam>
<lparam>Address:4177 16759</lparam>
<lparam>Address:4178 16760</lparam>
<lparam>Address:4179 16761</lparam>
<lparam>Address:4180 16768</lparam>
<lparam>Address:4181 16769</lparam>
<lparam>Address:4182 16770</lparam>
<lparam>Address:4183 16771</lparam>
<lparam>Address:4184 16772</lparam>
<lparam>Address:4185 16773</lparam>
<lparam>Address:4186 16774</lparam>
<lparam>Address:4187 16775</lparam>
<lparam>Address:4188 16776</lparam>
<lparam>Address:4189 16777</lparam>
<lparam>Address:4190 16784</lparam>
<lparam>Address:4191 16785</lparam>
<lparam>Address:4192 16786</lparam>
<lparam>Address:4193 16787</lparam>
<lparam>Address:4194 16788</lparam>
<lparam>Address:4195 16789</lparam>
<lparam>Address:4196 16790</lparam>
<lparam>Address:4197 16791</lparam>
<lparam>Address:4198 16792</lparam>
<lparam>Address:4199 16793</lparam>
<lparam>Address:4200 16896</lparam>
<lparam>Address:4201 16897</lparam>
<lparam>Address:4202 16898</lparam>
<lparam>Address:4203 16899</lparam>
<lparam>Address:4204 16900</lparam>
<lparam>Address:4205 16901</lparam>
<lparam>Address:4206 16902</lparam>
<lparam>Address:4207 16903</lparam>
<lparam>Address:4208 16904</lparam>
<lparam>Address:4209 16905</lparam>
<lparam>Address:4210 16912</lparam>
<lparam>Address:4211 16913</lparam>
<lparam>Address:4212 16914</lparam>
<lparam>Address:4213 16915</lparam>
<lparam>Address:4214 16916</lparam>
<lparam>Address:4215 16917</lparam>
<lparam>Address:4216 16918</lparam>
<lparam>Address:4217 16919</lparam>
<lparam>Address:4218 16920</lparam>
<lparam>Address:4219 16921</lparam>
<lparam>Address:4220 16928</lparam>
<lparam>Address:4221 16929</lparam>
<lparam>Address:4222 16930</lparam>
<lparam>Address:4223 16931</lparam>
<lparam>Address:4224 16932</lparam>
<lparam>Address:4225 16933</lparam>
<lparam>Address:4226 16934</lparam>
<lparam>Address:4227 16935</lparam>
<lparam>Address:4228 16936</lparam>
<lparam>Address:4229 16937</lparam>
<lparam>Address:4230 16944</lparam>
<lparam>Address:4231 16945</lparam>
<lparam>Address:4232 16946</lparam>
<lparam>Address:4233 16947</lparam>
<lparam>Address:4234 16948</lparam>
<lparam>Address:4235 16949</lparam>
<lparam>Address:4236 16950</lparam>
<lparam>Address:4237 16951</lparam>
<lparam>Address:4238 16952</lparam>
<lparam>Address:4239 16953</lparam>
<lparam>Address:4240 16960</lparam>
<lparam>Address:4241 16961</lparam>
<lparam>Address:4242 16962</lparam>
<lparam>Address:4243 16963</lparam>
<lparam>Address:4244 16964</lparam>
<lparam>Address:4245 16965</lparam>
<lparam>Address:4246 16966</lparam>
<lparam>Address:4247 16967</lparam>
<lparam>Address:4248 16968</lparam>
<lparam>Address:4249 16969</lparam>
<lparam>Address:4250 16976</lparam>
<lparam>Address:4251 16977</lparam>
<lparam>Address:4252 16978</lparam>
<lparam>Address:4253 16979</lparam>
<lparam>Address:4254 16980</lparam>
<lparam>Address:4255 16981</lparam>
<lparam>Address:4256 16982</lparam>
<lparam>Address:4257 16983</lparam>
<lparam>Address:4258 16984</lparam>
<lparam>Address:4259 16985</lparam>
<lparam>Address:4260 16992</lparam>
<lparam>Address:4261 16993</lparam>
<lparam>Address:4262 16994</lparam>
<lparam>Address:4263 16995</lparam>
<lparam>Address:4264 16996</lparam>
<lparam>Address:4265 16997</lparam>
<lparam>Address:4266 16998</lparam>
<lparam>Address:4267 16999</lparam>
<lparam>Address:4268 17000</lparam>
<lparam>Address:4269 17001</lparam>
<lparam>Address:4270 17008</lparam>
<lparam>Address:4271 17009</lparam>
<lparam>Address:4272 17010</lparam>
<lparam>Address:4273 17011</lparam>
<lparam>Address:4274 17012</lparam>
<lparam>Address:4275 17013</lparam>
<lparam>Address:4276 17014</lparam>
<lparam>Address:4277 17015</lparam>
<lparam>Address:4278 17016</lparam>
<lparam>Address:4279 17017</lparam>
<lparam>Address:4280 17024</lparam>
<lparam>Address:4281 17025</lparam>
<lparam>Address:4282 17026</lparam>
<lparam>Address:4283 17027</lparam>
<lparam>Address:4284 17028</lparam>
<lparam>Address:4285 17029</lparam>
<lparam>Address:4286 17030</lparam>
<lparam>Address:4287 17031</lparam>
<lparam>Address:4288 17032</lparam>
<lparam>Address:4289 17033</lparam>
<lparam>Address:4290 17040</lparam>
<lparam>Address:4291 17041</lparam>
<lparam>Address:4292 17042</lparam>
<lparam>Address:4293 17043</lparam>
<lparam>Address:4294 17044</lparam>
<lparam>Address:4295 17045</lparam>
<lparam>Address:4296 17046</lparam>
<lparam>Address:4297 17047</lparam>
<lparam>Address:4298 17048</lparam>
<lparam>Address:4299 17049</lparam>
<lparam>Address:4300 17152</lparam>
<lparam>Address:4301 17153</lparam>
<lparam>Address:4302 17154</lparam>
<lparam>Address:4303 17155</lparam>
<lparam>Address:4304 17156</lparam>
<lparam>Address:4305 17157</lparam>
<lparam>Address:4306 17158</lparam>
<lparam>Address:4307 17159</lparam>
<lparam>Address:4308 17160</lparam>
<lparam>Address:4309 17161</lparam>
<lparam>Address:4310 17168</lparam>
<lparam>Address:4311 17169</lparam>
<lparam>Address:4312 17170</lparam>
<lparam>Address:4313 17171</lparam>
<lparam>Address:4314 17172</lparam>
<lparam>Address:4315 17173</lparam>
<lparam>Address:4316 17174</lparam>
<lparam>Address:4317 17175</lparam>
<lparam>Address:4318 17176</lparam>
<lparam>Address:4319 17177</lparam>
<lparam>Address:4320 17184</lparam>
<lparam>Address:4321 17185</lparam>
<lparam>Address:4322 17186</lparam>
<lparam>Address:4323 17187</lparam>
<lparam>Address:4324 17188</lparam>
<lparam>Address:4325 17189</lparam>
<lparam>Address:4326 17190</lparam>
<lparam>Address:4327 17191</lparam>
<lparam>Address:4328 17192</lparam>
<lparam>Address:4329 17193</lparam>
<lparam>Address:4330 17200</lparam>
<lparam>Address:4331 17201</lparam>
<lparam>Address:4332 17202</lparam>
<lparam>Address:4333 17203</lparam>
<lparam>Address:4334 17204</lparam>
<lparam>Address:4335 17205</lparam>
<lparam>Address:4336 17206</lparam>
<lparam>Address:4337 17207</lparam>
<lparam>Address:4338 17208</lparam>
<lparam>Address:4339 17209</lparam>
<lparam>Address:4340 17216</lparam>
<lparam>Address:4341 17217</lparam>
<lparam>Address:4342 17218</lparam>
<lparam>Address:4343 17219</lparam>
<lparam>Address:4344 17220</lparam>
<lparam>Address:4345 17221</lparam>
<lparam>Address:4346 17222</lparam>
<lparam>Address:4347 17223</lparam>
<lparam>Address:4348 17224</lparam>
<lparam>Address:4349 17225</lparam>
<lparam>Address:4350 17232</lparam>
<lparam>Address:4351 17233</lparam>
<lparam>Address:4352 17234</lparam>
<lparam>Address:4353 17235</lparam>
<lparam>Address:4354 17236</lparam>
<lparam>Address:4355 17237</lparam>
<lparam>Address:4356 17238</lparam>
<lparam>Address:4357 17239</lparam>
<lparam>Address:4358 17240</lparam>
<lparam>Address:4359 17241</lparam>
<lparam>Address:4360 17248</lparam>
<lparam>Address:4361 17249</lparam>
<lparam>Address:4362 17250</lparam>
<lparam>Address:4363 17251</lparam>
<lparam>Address:4364 17252</lparam>
<lparam>Address:4365 17253</lparam>
<lparam>Address:4366 17254</lparam>
<lparam>Address:4367 17255</lparam>
<lparam>Address:4368 17256</lparam>
<lparam>Address:4369 17257</lparam>
<lparam>Address:4370 17264</lparam>
<lparam>Address:4371 17265</lparam>
<lparam>Address:4372 17266</lparam>
<lparam>Address:4373 17267</lparam>
<lparam>Address:4374 17268</lparam>
<lparam>Address:4375 17269</lparam>
<lparam>Address:4376 17270</lparam>
<lparam>Address:4377 17271</lparam>
<lparam>Address:4378 17272</lparam>
<lparam>Address:4379 17273</lparam>
<lparam>Address:4380 17280</lparam>
<lparam>Address:4381 17281</lparam>
<lparam>Address:4382 17282</lparam>
<lparam>Address:4383 17283</lparam>
<lparam>Address:4384 17284</lparam>
<lparam>Address:4385 17285</lparam>
<lparam>Address:4386 17286</lparam>
<lparam>Address:4387 17287</lparam>
<lparam>Address:4388 17288</lparam>
<lparam>Address:4389 17289</lparam>
<lparam>Address:4390 17296</lparam>
<lparam>Address:4391 17297</lparam>
<lparam>Address:4392 17298</lparam>
<lparam>Address:4393 17299</lparam>
<lparam>Address:4394 17300</lparam>
<lparam>Address:4395 17301</lparam>
<lparam>Address:4396 17302</lparam>
<lparam>Address:4397 17303</lparam>
<lparam>Address:4398 17304</lparam>
<lparam>Address:4399 17305</lparam>
<lparam>Address:4400 17408</lparam>
<lparam>Address:4401 17409</lparam>
<lparam>Address:4402 17410</lparam>
<lparam>Address:4403 17411</lparam>
<lparam>Address:4404 17412</lparam>
<lparam>Address:4405 17413</lparam>
<lparam>Address:4406 17414</lparam>
<lparam>Address:4407 17415</lparam>
<lparam>Address:4408 17416</lparam>
<lparam>Address:4409 17417</lparam>
<lparam>Address:4410 17424</lparam>
<lparam>Address:4411 17425</lparam>
<lparam>Address:4412 17426</lparam>
<lparam>Address:4413 17427</lparam>
<lparam>Address:4414 17428</lparam>
<lparam>Address:4415 17429</lparam>
<lparam>Address:4416 17430</lparam>
<lparam>Address:4417 17431</lparam>
<lparam>Address:4418 17432</lparam>
<lparam>Address:4419 17433</lparam>
<lparam>Address:4420 17440</lparam>
<lparam>Address:4421 17441</lparam>
<lparam>Address:4422 17442</lparam>
<lparam>Address:4423 17443</lparam>
<lparam>Address:4424 17444</lparam>
<lparam>Address:4425 17445</lparam>
<lparam>Address:4426 17446</lparam>
<lparam>Address:4427 17447</lparam>
<lparam>Address:4428 17448</lparam>
<lparam>Address:4429 17449</lparam>
<lparam>Address:4430 17456</lparam>
<lparam>Address:4431 17457</lparam>
<lparam>Address:4432 17458</lparam>
<lparam>Address:4433 17459</lparam>
<lparam>Address:4434 17460</lparam>
<lparam>Address:4435 17461</lparam>
<lparam>Address:4436 17462</lparam>
<lparam>Address:4437 17463</lparam>
<lparam>Address:4438 17464</lparam>
<lparam>Address:4439 17465</lparam>
<lparam>Address:4440 17472</lparam>
<lparam>Address:4441 17473</lparam>
<lparam>Address:4442 17474</lparam>
<lparam>Address:4443 17475</lparam>
<lparam>Address:4444 17476</lparam>
<lparam>Address:4445 17477</lparam>
<lparam>Address:4446 17478</lparam>
<lparam>Address:4447 17479</lparam>
<lparam>Address:4448 17480</lparam>
<lparam>Address:4449 17481</lparam>
<lparam>Address:4450 17488</lparam>
<lparam>Address:4451 17489</lparam>
<lparam>Address:4452 17490</lparam>
<lparam>Address:4453 17491</lparam>
<lparam>Address:4454 17492</lparam>
<lparam>Address:4455 17493</lparam>
<lparam>Address:4456 17494</lparam>
<lparam>Address:4457 17495</lparam>
<lparam>Address:4458 17496</lparam>
<lparam>Address:4459 17497</lparam>
<lparam>Address:4460 17504</lparam>
<lparam>Address:4461 17505</lparam>
<lparam>Address:4462 17506</lparam>
<lparam>Address:4463 17507</lparam>
<lparam>Address:4464 17508</lparam>
<lparam>Address:4465 17509</lparam>
<lparam>Address:4466 17510</lparam>
<lparam>Address:4467 17511</lparam>
<lparam>Address:4468 17512</lparam>
<lparam>Address:4469 17513</lparam>
<lparam>Address:4470 17520</lparam>
<lparam>Address:4471 17521</lparam>
<lparam>Address:4472 17522</lparam>
<lparam>Address:4473 17523</lparam>
<lparam>Address:4474 17524</lparam>
<lparam>Address:4475 17525</lparam>
<lparam>Address:4476 17526</lparam>
<lparam>Address:4477 17527</lparam>
<lparam>Address:4478 17528</lparam>
<lparam>Address:4479 17529</lparam>
<lparam>Address:4480 17536</lparam>
<lparam>Address:4481 17537</lparam>
<lparam>Address:4482 17538</lparam>
<lparam>Address:4483 17539</lparam>
<lparam>Address:4484 17540</lparam>
<lparam>Address:4485 17541</lparam>
<lparam>Address:4486 17542</lparam>
<lparam>Address:4487 17543</lparam>
<lparam>Address:4488 17544</lparam>
<lparam>Address:4489 17545</lparam>
<lparam>Address:4490 17552</lparam>
<lparam>Address:4491 17553</lparam>
<lparam>Address:4492 17554</lparam>
<lparam>Address:4493 17555</lparam>
<lparam>Address:4494 17556</lparam>
<lparam>Address:4495 17557</lparam>
<lparam>Address:4496 17558</lparam>
<lparam>Address:4497 17559</lparam>
<lparam>Address:4498 17560</lparam>
<lparam>Address:4499 17561</lparam>
<lparam>Address:4500 17664</lparam>
<lparam>Address:4501 17665</lparam>
<lparam>Address:4502 17666</lparam>
<lparam>Address:4503 17667</lparam>
<lparam>Address:4504 17668</lparam>
<lparam>Address:4505 17669</lparam>
<lparam>Address:4506 17670</lparam>
<lparam>Address:4507 17671</lparam>
<lparam>Address:4508 17672</lparam>
<lparam>Address:4509 17673</lparam>
<lparam>Address:4510 17680</lparam>
<lparam>Address:4511 17681</lparam>
<lparam>Address:4512 17682</lparam>
<lparam>Address:4513 17683</lparam>
<lparam>Address:4514 17684</lparam>
<lparam>Address:4515 17685</lparam>
<lparam>Address:4516 17686</lparam>
<lparam>Address:4517 17687</lparam>
<lparam>Address:4518 17688</lparam>
<lparam>Address:4519 17689</lparam>
<lparam>Address:4520 17696</lparam>
<lparam>Address:4521 17697</lparam>
<lparam>Address:4522 17698</lparam>
<lparam>Address:4523 17699</lparam>
<lparam>Address:4524 17700</lparam>
<lparam>Address:4525 17701</lparam>
<lparam>Address:4526 17702</lparam>
<lparam>Address:4527 17703</lparam>
<lparam>Address:4528 17704</lparam>
<lparam>Address:4529 17705</lparam>
<lparam>Address:4530 17712</lparam>
<lparam>Address:4531 17713</lparam>
<lparam>Address:4532 17714</lparam>
<lparam>Address:4533 17715</lparam>
<lparam>Address:4534 17716</lparam>
<lparam>Address:4535 17717</lparam>
<lparam>Address:4536 17718</lparam>
<lparam>Address:4537 17719</lparam>
<lparam>Address:4538 17720</lparam>
<lparam>Address:4539 17721</lparam>
<lparam>Address:4540 17728</lparam>
<lparam>Address:4541 17729</lparam>
<lparam>Address:4542 17730</lparam>
<lparam>Address:4543 17731</lparam>
<lparam>Address:4544 17732</lparam>
<lparam>Address:4545 17733</lparam>
<lparam>Address:4546 17734</lparam>
<lparam>Address:4547 17735</lparam>
<lparam>Address:4548 17736</lparam>
<lparam>Address:4549 17737</lparam>
<lparam>Address:4550 17744</lparam>
<lparam>Address:4551 17745</lparam>
<lparam>Address:4552 17746</lparam>
<lparam>Address:4553 17747</lparam>
<lparam>Address:4554 17748</lparam>
<lparam>Address:4555 17749</lparam>
<lparam>Address:4556 17750</lparam>
<lparam>Address:4557 17751</lparam>
<lparam>Address:4558 17752</lparam>
<lparam>Address:4559 17753</lparam>
<lparam>Address:4560 17760</lparam>
<lparam>Address:4561 17761</lparam>
<lparam>Address:4562 17762</lparam>
<lparam>Address:4563 17763</lparam>
<lparam>Address:4564 17764</lparam>
<lparam>Address:4565 17765</lparam>
<lparam>Address:4566 17766</lparam>
<lparam>Address:4567 17767</lparam>
<lparam>Address:4568 17768</lparam>
<lparam>Address:4569 17769</lparam>
<lparam>Address:4570 17776</lparam>
<lparam>Address:4571 17777</lparam>
<lparam>Address:4572 17778</lparam>
<lparam>Address:4573 17779</lparam>
<lparam>Address:4574 17780</lparam>
<lparam>Address:4575 17781</lparam>
<lparam>Address:4576 17782</lparam>
<lparam>Address:4577 17783</lparam>
<lparam>Address:4578 17784</lparam>
<lparam>Address:4579 17785</lparam>
<lparam>Address:4580 17792</lparam>
<lparam>Address:4581 17793</lparam>
<lparam>Address:4582 17794</lparam>
<lparam>Address:4583 17795</lparam>
<lparam>Address:4584 17796</lparam>
<lparam>Address:4585 17797</lparam>
<lparam>Address:4586 17798</lparam>
<lparam>Address:4587 17799</lparam>
<lparam>Address:4588 17800</lparam>
<lparam>Address:4589 17801</lparam>
<lparam>Address:4590 17808</lparam>
<lparam>Address:4591 17809</lparam>
<lparam>Address:4592 17810</lparam>
<lparam>Address:4593 17811</lparam>
<lparam>Address:4594 17812</lparam>
<lparam>Address:4595 17813</lparam>
<lparam>Address:4596 17814</lparam>
<lparam>Address:4597 17815</lparam>
<lparam>Address:4598 17816</lparam>
<lparam>Address:4599 17817</lparam>
<lparam>Address:4600 17920</lparam>
<lparam>Address:4601 17921</lparam>
<lparam>Address:4602 17922</lparam>
<lparam>Address:4603 17923</lparam>
<lparam>Address:4604 17924</lparam>
<lparam>Address:4605 17925</lparam>
<lparam>Address:4606 17926</lparam>
<lparam>Address:4607 17927</lparam>
<lparam>Address:4608 17928</lparam>
<lparam>Address:4609 17929</lparam>
<lparam>Address:4610 17936</lparam>
<lparam>Address:4611 17937</lparam>
<lparam>Address:4612 17938</lparam>
<lparam>Address:4613 17939</lparam>
<lparam>Address:4614 17940</lparam>
<lparam>Address:4615 17941</lparam>
<lparam>Address:4616 17942</lparam>
<lparam>Address:4617 17943</lparam>
<lparam>Address:4618 17944</lparam>
<lparam>Address:4619 17945</lparam>
<lparam>Address:4620 17952</lparam>
<lparam>Address:4621 17953</lparam>
<lparam>Address:4622 17954</lparam>
<lparam>Address:4623 17955</lparam>
<lparam>Address:4624 17956</lparam>
<lparam>Address:4625 17957</lparam>
<lparam>Address:4626 17958</lparam>
<lparam>Address:4627 17959</lparam>
<lparam>Address:4628 17960</lparam>
<lparam>Address:4629 17961</lparam>
<lparam>Address:4630 17968</lparam>
<lparam>Address:4631 17969</lparam>
<lparam>Address:4632 17970</lparam>
<lparam>Address:4633 17971</lparam>
<lparam>Address:4634 17972</lparam>
<lparam>Address:4635 17973</lparam>
<lparam>Address:4636 17974</lparam>
<lparam>Address:4637 17975</lparam>
<lparam>Address:4638 17976</lparam>
<lparam>Address:4639 17977</lparam>
<lparam>Address:4640 17984</lparam>
<lparam>Address:4641 17985</lparam>
<lparam>Address:4642 17986</lparam>
<lparam>Address:4643 17987</lparam>
<lparam>Address:4644 17988</lparam>
<lparam>Address:4645 17989</lparam>
<lparam>Address:4646 17990</lparam>
<lparam>Address:4647 17991</lparam>
<lparam>Address:4648 17992</lparam>
<lparam>Address:4649 17993</lparam>
<lparam>Address:4650 18000</lparam>
<lparam>Address:4651 18001</lparam>
<lparam>Address:4652 18002</lparam>
<lparam>Address:4653 18003</lparam>
<lparam>Address:4654 18004</lparam>
<lparam>Address:4655 18005</lparam>
<lparam>Address:4656 18006</lparam>
<lparam>Address:4657 18007</lparam>
<lparam>Address:4658 18008</lparam>
<lparam>Address:4659 18009</lparam>
<lparam>Address:4660 18016</lparam>
<lparam>Address:4661 18017</lparam>
<lparam>Address:4662 18018</lparam>
<lparam>Address:4663 18019</lparam>
<lparam>Address:4664 18020</lparam>
<lparam>Address:4665 18021</lparam>
<lparam>Address:4666 18022</lparam>
<lparam>Address:4667 18023</lparam>
<lparam>Address:4668 18024</lparam>
<lparam>Address:4669 18025</lparam>
<lparam>Address:4670 18032</lparam>
<lparam>Address:4671 18033</lparam>
<lparam>Address:4672 18034</lparam>
<lparam>Address:4673 18035</lparam>
<lparam>Address:4674 18036</lparam>
<lparam>Address:4675 18037</lparam>
<lparam>Address:4676 18038</lparam>
<lparam>Address:4677 18039</lparam>
<lparam>Address:4678 18040</lparam>
<lparam>Address:4679 18041</lparam>
<lparam>Address:4680 18048</lparam>
<lparam>Address:4681 18049</lparam>
<lparam>Address:4682 18050</lparam>
<lparam>Address:4683 18051</lparam>
<lparam>Address:4684 18052</lparam>
<lparam>Address:4685 18053</lparam>
<lparam>Address:4686 18054</lparam>
<lparam>Address:4687 18055</lparam>
<lparam>Address:4688 18056</lparam>
<lparam>Address:4689 18057</lparam>
<lparam>Address:4690 18064</lparam>
<lparam>Address:4691 18065</lparam>
<lparam>Address:4692 18066</lparam>
<lparam>Address:4693 18067</lparam>
<lparam>Address:4694 18068</lparam>
<lparam>Address:4695 18069</lparam>
<lparam>Address:4696 18070</lparam>
<lparam>Address:4697 18071</lparam>
<lparam>Address:4698 18072</lparam>
<lparam>Address:4699 18073</lparam>
<lparam>Address:4700 18176</lparam>
<lparam>Address:4701 18177</lparam>
<lparam>Address:4702 18178</lparam>
<lparam>Address:4703 18179</lparam>
<lparam>Address:4704 18180</lparam>
<lparam>Address:4705 18181</lparam>
<lparam>Address:4706 18182</lparam>
<lparam>Address:4707 18183</lparam>
<lparam>Address:4708 18184</lparam>
<lparam>Address:4709 18185</lparam>
<lparam>Address:4710 18192</lparam>
<lparam>Address:4711 18193</lparam>
<lparam>Address:4712 18194</lparam>
<lparam>Address:4713 18195</lparam>
<lparam>Address:4714 18196</lparam>
<lparam>Address:4715 18197</lparam>
<lparam>Address:4716 18198</lparam>
<lparam>Address:4717 18199</lparam>
<lparam>Address:4718 18200</lparam>
<lparam>Address:4719 18201</lparam>
<lparam>Address:4720 18208</lparam>
<lparam>Address:4721 18209</lparam>
<lparam>Address:4722 18210</lparam>
<lparam>Address:4723 18211</lparam>
<lparam>Address:4724 18212</lparam>
<lparam>Address:4725 18213</lparam>
<lparam>Address:4726 18214</lparam>
<lparam>Address:4727 18215</lparam>
<lparam>Address:4728 18216</lparam>
<lparam>Address:4729 18217</lparam>
<lparam>Address:4730 18224</lparam>
<lparam>Address:4731 18225</lparam>
<lparam>Address:4732 18226</lparam>
<lparam>Address:4733 18227</lparam>
<lparam>Address:4734 18228</lparam>
<lparam>Address:4735 18229</lparam>
<lparam>Address:4736 18230</lparam>
<lparam>Address:4737 18231</lparam>
<lparam>Address:4738 18232</lparam>
<lparam>Address:4739 18233</lparam>
<lparam>Address:4740 18240</lparam>
<lparam>Address:4741 18241</lparam>
<lparam>Address:4742 18242</lparam>
<lparam>Address:4743 18243</lparam>
<lparam>Address:4744 18244</lparam>
<lparam>Address:4745 18245</lparam>
<lparam>Address:4746 18246</lparam>
<lparam>Address:4747 18247</lparam>
<lparam>Address:4748 18248</lparam>
<lparam>Address:4749 18249</lparam>
<lparam>Address:4750 18256</lparam>
<lparam>Address:4751 18257</lparam>
<lparam>Address:4752 18258</lparam>
<lparam>Address:4753 18259</lparam>
<lparam>Address:4754 18260</lparam>
<lparam>Address:4755 18261</lparam>
<lparam>Address:4756 18262</lparam>
<lparam>Address:4757 18263</lparam>
<lparam>Address:4758 18264</lparam>
<lparam>Address:4759 18265</lparam>
<lparam>Address:4760 18272</lparam>
<lparam>Address:4761 18273</lparam>
<lparam>Address:4762 18274</lparam>
<lparam>Address:4763 18275</lparam>
<lparam>Address:4764 18276</lparam>
<lparam>Address:4765 18277</lparam>
<lparam>Address:4766 18278</lparam>
<lparam>Address:4767 18279</lparam>
<lparam>Address:4768 18280</lparam>
<lparam>Address:4769 18281</lparam>
<lparam>Address:4770 18288</lparam>
<lparam>Address:4771 18289</lparam>
<lparam>Address:4772 18290</lparam>
<lparam>Address:4773 18291</lparam>
<lparam>Address:4774 18292</lparam>
<lparam>Address:4775 18293</lparam>
<lparam>Address:4776 18294</lparam>
<lparam>Address:4777 18295</lparam>
<lparam>Address:4778 18296</lparam>
<lparam>Address:4779 18297</lparam>
<lparam>Address:4780 18304</lparam>
<lparam>Address:4781 18305</lparam>
<lparam>Address:4782 18306</lparam>
<lparam>Address:4783 18307</lparam>
<lparam>Address:4784 18308</lparam>
<lparam>Address:4785 18309</lparam>
<lparam>Address:4786 18310</lparam>
<lparam>Address:4787 18311</lparam>
<lparam>Address:4788 18312</lparam>
<lparam>Address:4789 18313</lparam>
<lparam>Address:4790 18320</lparam>
<lparam>Address:4791 18321</lparam>
<lparam>Address:4792 18322</lparam>
<lparam>Address:4793 18323</lparam>
<lparam>Address:4794 18324</lparam>
<lparam>Address:4795 18325</lparam>
<lparam>Address:4796 18326</lparam>
<lparam>Address:4797 18327</lparam>
<lparam>Address:4798 18328</lparam>
<lparam>Address:4799 18329</lparam>
<lparam>Address:4800 18432</lparam>
<lparam>Address:4801 18433</lparam>
<lparam>Address:4802 18434</lparam>
<lparam>Address:4803 18435</lparam>
<lparam>Address:4804 18436</lparam>
<lparam>Address:4805 18437</lparam>
<lparam>Address:4806 18438</lparam>
<lparam>Address:4807 18439</lparam>
<lparam>Address:4808 18440</lparam>
<lparam>Address:4809 18441</lparam>
<lparam>Address:4810 18448</lparam>
<lparam>Address:4811 18449</lparam>
<lparam>Address:4812 18450</lparam>
<lparam>Address:4813 18451</lparam>
<lparam>Address:4814 18452</lparam>
<lparam>Address:4815 18453</lparam>
<lparam>Address:4816 18454</lparam>
<lparam>Address:4817 18455</lparam>
<lparam>Address:4818 18456</lparam>
<lparam>Address:4819 18457</lparam>
<lparam>Address:4820 18464</lparam>
<lparam>Address:4821 18465</lparam>
<lparam>Address:4822 18466</lparam>
<lparam>Address:4823 18467</lparam>
<lparam>Address:4824 18468</lparam>
<lparam>Address:4825 18469</lparam>
<lparam>Address:4826 18470</lparam>
<lparam>Address:4827 18471</lparam>
<lparam>Address:4828 18472</lparam>
<lparam>Address:4829 18473</lparam>
<lparam>Address:4830 18480</lparam>
<lparam>Address:4831 18481</lparam>
<lparam>Address:4832 18482</lparam>
<lparam>Address:4833 18483</lparam>
<lparam>Address:4834 18484</lparam>
<lparam>Address:4835 18485</lparam>
<lparam>Address:4836 18486</lparam>
<lparam>Address:4837 18487</lparam>
<lparam>Address:4838 18488</lparam>
<lparam>Address:4839 18489</lparam>
<lparam>Address:4840 18496</lparam>
<lparam>Address:4841 18497</lparam>
<lparam>Address:4842 18498</lparam>
<lparam>Address:4843 18499</lparam>
<lparam>Address:4844 18500</lparam>
<lparam>Address:4845 18501</lparam>
<lparam>Address:4846 18502</lparam>
<lparam>Address:4847 18503</lparam>
<lparam>Address:4848 18504</lparam>
<lparam>Address:4849 18505</lparam>
<lparam>Address:4850 18512</lparam>
<lparam>Address:4851 18513</lparam>
<lparam>Address:4852 18514</lparam>
<lparam>Address:4853 18515</lparam>
<lparam>Address:4854 18516</lparam>
<lparam>Address:4855 18517</lparam>
<lparam>Address:4856 18518</lparam>
<lparam>Address:4857 18519</lparam>
<lparam>Address:4858 18520</lparam>
<lparam>Address:4859 18521</lparam>
<lparam>Address:4860 18528</lparam>
<lparam>Address:4861 18529</lparam>
<lparam>Address:4862 18530</lparam>
<lparam>Address:4863 18531</lparam>
<lparam>Address:4864 18532</lparam>
<lparam>Address:4865 18533</lparam>
<lparam>Address:4866 18534</lparam>
<lparam>Address:4867 18535</lparam>
<lparam>Address:4868 18536</lparam>
<lparam>Address:4869 18537</lparam>
<lparam>Address:4870 18544</lparam>
<lparam>Address:4871 18545</lparam>
<lparam>Address:4872 18546</lparam>
<lparam>Address:4873 18547</lparam>
<lparam>Address:4874 18548</lparam>
<lparam>Address:4875 18549</lparam>
<lparam>Address:4876 18550</lparam>
<lparam>Address:4877 18551</lparam>
<lparam>Address:4878 18552</lparam>
<lparam>Address:4879 18553</lparam>
<lparam>Address:4880 18560</lparam>
<lparam>Address:4881 18561</lparam>
<lparam>Address:4882 18562</lparam>
<lparam>Address:4883 18563</lparam>
<lparam>Address:4884 18564</lparam>
<lparam>Address:4885 18565</lparam>
<lparam>Address:4886 18566</lparam>
<lparam>Address:4887 18567</lparam>
<lparam>Address:4888 18568</lparam>
<lparam>Address:4889 18569</lparam>
<lparam>Address:4890 18576</lparam>
<lparam>Address:4891 18577</lparam>
<lparam>Address:4892 18578</lparam>
<lparam>Address:4893 18579</lparam>
<lparam>Address:4894 18580</lparam>
<lparam>Address:4895 18581</lparam>
<lparam>Address:4896 18582</lparam>
<lparam>Address:4897 18583</lparam>
<lparam>Address:4898 18584</lparam>
<lparam>Address:4899 18585</lparam>
<lparam>Address:4900 18688</lparam>
<lparam>Address:4901 18689</lparam>
<lparam>Address:4902 18690</lparam>
<lparam>Address:4903 18691</lparam>
<lparam>Address:4904 18692</lparam>
<lparam>Address:4905 18693</lparam>
<lparam>Address:4906 18694</lparam>
<lparam>Address:4907 18695</lparam>
<lparam>Address:4908 18696</lparam>
<lparam>Address:4909 18697</lparam>
<lparam>Address:4910 18704</lparam>
<lparam>Address:4911 18705</lparam>
<lparam>Address:4912 18706</lparam>
<lparam>Address:4913 18707</lparam>
<lparam>Address:4914 18708</lparam>
<lparam>Address:4915 18709</lparam>
<lparam>Address:4916 18710</lparam>
<lparam>Address:4917 18711</lparam>
<lparam>Address:4918 18712</lparam>
<lparam>Address:4919 18713</lparam>
<lparam>Address:4920 18720</lparam>
<lparam>Address:4921 18721</lparam>
<lparam>Address:4922 18722</lparam>
<lparam>Address:4923 18723</lparam>
<lparam>Address:4924 18724</lparam>
<lparam>Address:4925 18725</lparam>
<lparam>Address:4926 18726</lparam>
<lparam>Address:4927 18727</lparam>
<lparam>Address:4928 18728</lparam>
<lparam>Address:4929 18729</lparam>
<lparam>Address:4930 18736</lparam>
<lparam>Address:4931 18737</lparam>
<lparam>Address:4932 18738</lparam>
<lparam>Address:4933 18739</lparam>
<lparam>Address:4934 18740</lparam>
<lparam>Address:4935 18741</lparam>
<lparam>Address:4936 18742</lparam>
<lparam>Address:4937 18743</lparam>
<lparam>Address:4938 18744</lparam>
<lparam>Address:4939 18745</lparam>
<lparam>Address:4940 18752</lparam>
<lparam>Address:4941 18753</lparam>
<lparam>Address:4942 18754</lparam>
<lparam>Address:4943 18755</lparam>
<lparam>Address:4944 18756</lparam>
<lparam>Address:4945 18757</lparam>
<lparam>Address:4946 18758</lparam>
<lparam>Address:4947 18759</lparam>
<lparam>Address:4948 18760</lparam>
<lparam>Address:4949 18761</lparam>
<lparam>Address:4950 18768</lparam>
<lparam>Address:4951 18769</lparam>
<lparam>Address:4952 18770</lparam>
<lparam>Address:4953 18771</lparam>
<lparam>Address:4954 18772</lparam>
<lparam>Address:4955 18773</lparam>
<lparam>Address:4956 18774</lparam>
<lparam>Address:4957 18775</lparam>
<lparam>Address:4958 18776</lparam>
<lparam>Address:4959 18777</lparam>
<lparam>Address:4960 18784</lparam>
<lparam>Address:4961 18785</lparam>
<lparam>Address:4962 18786</lparam>
<lparam>Address:4963 18787</lparam>
<lparam>Address:4964 18788</lparam>
<lparam>Address:4965 18789</lparam>
<lparam>Address:4966 18790</lparam>
<lparam>Address:4967 18791</lparam>
<lparam>Address:4968 18792</lparam>
<lparam>Address:4969 18793</lparam>
<lparam>Address:4970 18800</lparam>
<lparam>Address:4971 18801</lparam>
<lparam>Address:4972 18802</lparam>
<lparam>Address:4973 18803</lparam>
<lparam>Address:4974 18804</lparam>
<lparam>Address:4975 18805</lparam>
<lparam>Address:4976 18806</lparam>
<lparam>Address:4977 18807</lparam>
<lparam>Address:4978 18808</lparam>
<lparam>Address:4979 18809</lparam>
<lparam>Address:4980 18816</lparam>
<lparam>Address:4981 18817</lparam>
<lparam>Address:4982 18818</lparam>
<lparam>Address:4983 18819</lparam>
<lparam>Address:4984 18820</lparam>
<lparam>Address:4985 18821</lparam>
<lparam>Address:4986 18822</lparam>
<lparam>Address:4987 18823</lparam>
<lparam>Address:4988 18824</lparam>
<lparam>Address:4989 18825</lparam>
<lparam>Address:4990 18832</lparam>
<lparam>Address:4991 18833</lparam>
<lparam>Address:4992 18834</lparam>
<lparam>Address:4993 18835</lparam>
<lparam>Address:4994 18836</lparam>
<lparam>Address:4995 18837</lparam>
<lparam>Address:4996 18838</lparam>
<lparam>Address:4997 18839</lparam>
<lparam>Address:4998 18840</lparam>
<lparam>Address:4999 18841</lparam>
<lparam>Address:5000 16384</lparam>
<lparam>Address:5001 20481</lparam>
<lparam>Address:5002 20482</lparam>
<lparam>Address:5003 20483</lparam>
<lparam>Address:5004 20484</lparam>
<lparam>Address:5005 20485</lparam>
<lparam>Address:5006 20486</lparam>
<lparam>Address:5007 20487</lparam>
<lparam>Address:5008 20488</lparam>
<lparam>Address:5009 20489</lparam>
<lparam>Address:5010 20496</lparam>
<lparam>Address:5011 20497</lparam>
<lparam>Address:5012 20498</lparam>
<lparam>Address:5013 20499</lparam>
<lparam>Address:5014 20500</lparam>
<lparam>Address:5015 20501</lparam>
<lparam>Address:5016 20502</lparam>
<lparam>Address:5017 20503</lparam>
<lparam>Address:5018 20504</lparam>
<lparam>Address:5019 20505</lparam>
<lparam>Address:5020 20512</lparam>
<lparam>Address:5021 20513</lparam>
<lparam>Address:5022 20514</lparam>
<lparam>Address:5023 20515</lparam>
<lparam>Address:5024 20516</lparam>
<lparam>Address:5025 20517</lparam>
<lparam>Address:5026 20518</lparam>
<lparam>Address:5027 20519</lparam>
<lparam>Address:5028 20520</lparam>
<lparam>Address:5029 20521</lparam>
<lparam>Address:5030 20528</lparam>
<lparam>Address:5031 20529</lparam>
<lparam>Address:5032 20530</lparam>
<lparam>Address:5033 20531</lparam>
<lparam>Address:5034 20532</lparam>
<lparam>Address:5035 20533</lparam>
<lparam>Address:5036 20534</lparam>
<lparam>Address:5037 20535</lparam>
<lparam>Address:5038 20536</lparam>
<lparam>Address:5039 20537</lparam>
<lparam>Address:5040 20544</lparam>
<lparam>Address:5041 20545</lparam>
<lparam>Address:5042 20546</lparam>
<lparam>Address:5043 20547</lparam>
<lparam>Address:5044 20548</lparam>
<lparam>Address:5045 20549</lparam>
<lparam>Address:5046 20550</lparam>
<lparam>Address:5047 20551</lparam>
<lparam>Address:5048 20552</lparam>
<lparam>Address:5049 20553</lparam>
<lparam>Address:5050 20560</lparam>
<lparam>Address:5051 20561</lparam>
<lparam>Address:5052 20562</lparam>
<lparam>Address:5053 20563</lparam>
<lparam>Address:5054 20564</lparam>
<lparam>Address:5055 20565</lparam>
<lparam>Address:5056 20566</lparam>
<lparam>Address:5057 20567</lparam>
<lparam>Address:5058 20568</lparam>
<lparam>Address:5059 20569</lparam>
<lparam>Address:5060 20576</lparam>
<lparam>Address:5061 20577</lparam>
<lparam>Address:5062 20578</lparam>
<lparam>Address:5063 20579</lparam>
<lparam>Address:5064 20580</lparam>
<lparam>Address:5065 20581</lparam>
<lparam>Address:5066 20582</lparam>
<lparam>Address:5067 20583</lparam>
<lparam>Address:5068 20584</lparam>
<lparam>Address:5069 20585</lparam>
<lparam>Address:5070 20592</lparam>
<lparam>Address:5071 20593</lparam>
<lparam>Address:5072 20594</lparam>
<lparam>Address:5073 20595</lparam>
<lparam>Address:5074 20596</lparam>
<lparam>Address:5075 20597</lparam>
<lparam>Address:5076 20598</lparam>
<lparam>Address:5077 20599</lparam>
<lparam>Address:5078 20600</lparam>
<lparam>Address:5079 20601</lparam>
<lparam>Address:5080 20608</lparam>
<lparam>Address:5081 20609</lparam>
<lparam>Address:5082 20610</lparam>
<lparam>Address:5083 20611</lparam>
<lparam>Address:5084 20612</lparam>
<lparam>Address:5085 20613</lparam>
<lparam>Address:5086 20614</lparam>
<lparam>Address:5087 20615</lparam>
<lparam>Address:5088 20616</lparam>
<lparam>Address:5089 20617</lparam>
<lparam>Address:5090 20624</lparam>
<lparam>Address:5091 20625</lparam>
<lparam>Address:5092 20626</lparam>
<lparam>Address:5093 20627</lparam>
<lparam>Address:5094 20628</lparam>
<lparam>Address:5095 20629</lparam>
<lparam>Address:5096 20630</lparam>
<lparam>Address:5097 20631</lparam>
<lparam>Address:5098 20632</lparam>
<lparam>Address:5099 20633</lparam>
<lparam>Address:5100 20736</lparam>
<lparam>Address:5101 20737</lparam>
<lparam>Address:5102 20738</lparam>
<lparam>Address:5103 20739</lparam>
<lparam>Address:5104 20740</lparam>
<lparam>Address:5105 20741</lparam>
<lparam>Address:5106 20742</lparam>
<lparam>Address:5107 20743</lparam>
<lparam>Address:5108 20744</lparam>
<lparam>Address:5109 20745</lparam>
<lparam>Address:5110 20752</lparam>
<lparam>Address:5111 20753</lparam>
<lparam>Address:5112 20754</lparam>
<lparam>Address:5113 20755</lparam>
<lparam>Address:5114 20756</lparam>
<lparam>Address:5115 20757</lparam>
<lparam>Address:5116 20758</lparam>
<lparam>Address:5117 20759</lparam>
<lparam>Address:5118 20760</lparam>
<lparam>Address:5119 20761</lparam>
<lparam>Address:5120 20768</lparam>
<lparam>Address:5121 20769</lparam>
<lparam>Address:5122 20770</lparam>
<lparam>Address:5123 20771</lparam>
<lparam>Address:5124 20772</lparam>
<lparam>Address:5125 20773</lparam>
<lparam>Address:5126 20774</lparam>
<lparam>Address:5127 20775</lparam>
<lparam>Address:5128 20776</lparam>
<lparam>Address:5129 20777</lparam>
<lparam>Address:5130 20784</lparam>
<lparam>Address:5131 20785</lparam>
<lparam>Address:5132 20786</lparam>
<lparam>Address:5133 20787</lparam>
<lparam>Address:5134 20788</lparam>
<lparam>Address:5135 20789</lparam>
<lparam>Address:5136 20790</lparam>
<lparam>Address:5137 20791</lparam>
<lparam>Address:5138 20792</lparam>
<lparam>Address:5139 20793</lparam>
<lparam>Address:5140 20800</lparam>
<lparam>Address:5141 20801</lparam>
<lparam>Address:5142 20802</lparam>
<lparam>Address:5143 20803</lparam>
<lparam>Address:5144 20804</lparam>
<lparam>Address:5145 20805</lparam>
<lparam>Address:5146 20806</lparam>
<lparam>Address:5147 20807</lparam>
<lparam>Address:5148 20808</lparam>
<lparam>Address:5149 20809</lparam>
<lparam>Address:5150 20816</lparam>
<lparam>Address:5151 20817</lparam>
<lparam>Address:5152 20818</lparam>
<lparam>Address:5153 20819</lparam>
<lparam>Address:5154 20820</lparam>
<lparam>Address:5155 20821</lparam>
<lparam>Address:5156 20822</lparam>
<lparam>Address:5157 20823</lparam>
<lparam>Address:5158 20824</lparam>
<lparam>Address:5159 20825</lparam>
<lparam>Address:5160 20832</lparam>
<lparam>Address:5161 20833</lparam>
<lparam>Address:5162 20834</lparam>
<lparam>Address:5163 20835</lparam>
<lparam>Address:5164 20836</lparam>
<lparam>Address:5165 20837</lparam>
<lparam>Address:5166 20838</lparam>
<lparam>Address:5167 20839</lparam>
<lparam>Address:5168 20840</lparam>
<lparam>Address:5169 20841</lparam>
<lparam>Address:5170 20848</lparam>
<lparam>Address:5171 20849</lparam>
<lparam>Address:5172 20850</lparam>
<lparam>Address:5173 20851</lparam>
<lparam>Address:5174 20852</lparam>
<lparam>Address:5175 20853</lparam>
<lparam>Address:5176 20854</lparam>
<lparam>Address:5177 20855</lparam>
<lparam>Address:5178 20856</lparam>
<lparam>Address:5179 20857</lparam>
<lparam>Address:5180 20864</lparam>
<lparam>Address:5181 20865</lparam>
<lparam>Address:5182 20866</lparam>
<lparam>Address:5183 20867</lparam>
<lparam>Address:5184 20868</lparam>
<lparam>Address:5185 20869</lparam>
<lparam>Address:5186 20870</lparam>
<lparam>Address:5187 20871</lparam>
<lparam>Address:5188 20872</lparam>
<lparam>Address:5189 20873</lparam>
<lparam>Address:5190 20880</lparam>
<lparam>Address:5191 20881</lparam>
<lparam>Address:5192 20882</lparam>
<lparam>Address:5193 20883</lparam>
<lparam>Address:5194 20884</lparam>
<lparam>Address:5195 20885</lparam>
<lparam>Address:5196 20886</lparam>
<lparam>Address:5197 20887</lparam>
<lparam>Address:5198 20888</lparam>
<lparam>Address:5199 20889</lparam>
<lparam>Address:5200 20992</lparam>
<lparam>Address:5201 20993</lparam>
<lparam>Address:5202 20994</lparam>
<lparam>Address:5203 20995</lparam>
<lparam>Address:5204 20996</lparam>
<lparam>Address:5205 20997</lparam>
<lparam>Address:5206 20998</lparam>
<lparam>Address:5207 20999</lparam>
<lparam>Address:5208 21000</lparam>
<lparam>Address:5209 21001</lparam>
<lparam>Address:5210 21008</lparam>
<lparam>Address:5211 21009</lparam>
<lparam>Address:5212 21010</lparam>
<lparam>Address:5213 21011</lparam>
<lparam>Address:5214 21012</lparam>
<lparam>Address:5215 21013</lparam>
<lparam>Address:5216 21014</lparam>
<lparam>Address:5217 21015</lparam>
<lparam>Address:5218 21016</lparam>
<lparam>Address:5219 21017</lparam>
<lparam>Address:5220 21024</lparam>
<lparam>Address:5221 21025</lparam>
<lparam>Address:5222 21026</lparam>
<lparam>Address:5223 21027</lparam>
<lparam>Address:5224 21028</lparam>
<lparam>Address:5225 21029</lparam>
<lparam>Address:5226 21030</lparam>
<lparam>Address:5227 21031</lparam>
<lparam>Address:5228 21032</lparam>
<lparam>Address:5229 21033</lparam>
<lparam>Address:5230 21040</lparam>
<lparam>Address:5231 21041</lparam>
<lparam>Address:5232 21042</lparam>
<lparam>Address:5233 21043</lparam>
<lparam>Address:5234 21044</lparam>
<lparam>Address:5235 21045</lparam>
<lparam>Address:5236 21046</lparam>
<lparam>Address:5237 21047</lparam>
<lparam>Address:5238 21048</lparam>
<lparam>Address:5239 21049</lparam>
<lparam>Address:5240 21056</lparam>
<lparam>Address:5241 21057</lparam>
<lparam>Address:5242 21058</lparam>
<lparam>Address:5243 21059</lparam>
<lparam>Address:5244 21060</lparam>
<lparam>Address:5245 21061</lparam>
<lparam>Address:5246 21062</lparam>
<lparam>Address:5247 21063</lparam>
<lparam>Address:5248 21064</lparam>
<lparam>Address:5249 21065</lparam>
<lparam>Address:5250 21072</lparam>
<lparam>Address:5251 21073</lparam>
<lparam>Address:5252 21074</lparam>
<lparam>Address:5253 21075</lparam>
<lparam>Address:5254 21076</lparam>
<lparam>Address:5255 21077</lparam>
<lparam>Address:5256 21078</lparam>
<lparam>Address:5257 21079</lparam>
<lparam>Address:5258 21080</lparam>
<lparam>Address:5259 21081</lparam>
<lparam>Address:5260 21088</lparam>
<lparam>Address:5261 21089</lparam>
<lparam>Address:5262 21090</lparam>
<lparam>Address:5263 21091</lparam>
<lparam>Address:5264 21092</lparam>
<lparam>Address:5265 21093</lparam>
<lparam>Address:5266 21094</lparam>
<lparam>Address:5267 21095</lparam>
<lparam>Address:5268 21096</lparam>
<lparam>Address:5269 21097</lparam>
<lparam>Address:5270 21104</lparam>
<lparam>Address:5271 21105</lparam>
<lparam>Address:5272 21106</lparam>
<lparam>Address:5273 21107</lparam>
<lparam>Address:5274 21108</lparam>
<lparam>Address:5275 21109</lparam>
<lparam>Address:5276 21110</lparam>
<lparam>Address:5277 21111</lparam>
<lparam>Address:5278 21112</lparam>
<lparam>Address:5279 21113</lparam>
<lparam>Address:5280 21120</lparam>
<lparam>Address:5281 21121</lparam>
<lparam>Address:5282 21122</lparam>
<lparam>Address:5283 21123</lparam>
<lparam>Address:5284 21124</lparam>
<lparam>Address:5285 21125</lparam>
<lparam>Address:5286 21126</lparam>
<lparam>Address:5287 21127</lparam>
<lparam>Address:5288 21128</lparam>
<lparam>Address:5289 21129</lparam>
<lparam>Address:5290 21136</lparam>
<lparam>Address:5291 21137</lparam>
<lparam>Address:5292 21138</lparam>
<lparam>Address:5293 21139</lparam>
<lparam>Address:5294 21140</lparam>
<lparam>Address:5295 21141</lparam>
<lparam>Address:5296 21142</lparam>
<lparam>Address:5297 21143</lparam>
<lparam>Address:5298 21144</lparam>
<lparam>Address:5299 21145</lparam>
<lparam>Address:5300 21248</lparam>
<lparam>Address:5301 21249</lparam>
<lparam>Address:5302 21250</lparam>
<lparam>Address:5303 21251</lparam>
<lparam>Address:5304 21252</lparam>
<lparam>Address:5305 21253</lparam>
<lparam>Address:5306 21254</lparam>
<lparam>Address:5307 21255</lparam>
<lparam>Address:5308 21256</lparam>
<lparam>Address:5309 21257</lparam>
<lparam>Address:5310 21264</lparam>
<lparam>Address:5311 21265</lparam>
<lparam>Address:5312 21266</lparam>
<lparam>Address:5313 21267</lparam>
<lparam>Address:5314 21268</lparam>
<lparam>Address:5315 21269</lparam>
<lparam>Address:5316 21270</lparam>
<lparam>Address:5317 21271</lparam>
<lparam>Address:5318 21272</lparam>
<lparam>Address:5319 21273</lparam>
<lparam>Address:5320 21280</lparam>
<lparam>Address:5321 21281</lparam>
<lparam>Address:5322 21282</lparam>
<lparam>Address:5323 21283</lparam>
<lparam>Address:5324 21284</lparam>
<lparam>Address:5325 21285</lparam>
<lparam>Address:5326 21286</lparam>
<lparam>Address:5327 21287</lparam>
<lparam>Address:5328 21288</lparam>
<lparam>Address:5329 21289</lparam>
<lparam>Address:5330 21296</lparam>
<lparam>Address:5331 21297</lparam>
<lparam>Address:5332 21298</lparam>
<lparam>Address:5333 21299</lparam>
<lparam>Address:5334 21300</lparam>
<lparam>Address:5335 21301</lparam>
<lparam>Address:5336 21302</lparam>
<lparam>Address:5337 21303</lparam>
<lparam>Address:5338 21304</lparam>
<lparam>Address:5339 21305</lparam>
<lparam>Address:5340 21312</lparam>
<lparam>Address:5341 21313</lparam>
<lparam>Address:5342 21314</lparam>
<lparam>Address:5343 21315</lparam>
<lparam>Address:5344 21316</lparam>
<lparam>Address:5345 21317</lparam>
<lparam>Address:5346 21318</lparam>
<lparam>Address:5347 21319</lparam>
<lparam>Address:5348 21320</lparam>
<lparam>Address:5349 21321</lparam>
<lparam>Address:5350 21328</lparam>
<lparam>Address:5351 21329</lparam>
<lparam>Address:5352 21330</lparam>
<lparam>Address:5353 21331</lparam>
<lparam>Address:5354 21332</lparam>
<lparam>Address:5355 21333</lparam>
<lparam>Address:5356 21334</lparam>
<lparam>Address:5357 21335</lparam>
<lparam>Address:5358 21336</lparam>
<lparam>Address:5359 21337</lparam>
<lparam>Address:5360 21344</lparam>
<lparam>Address:5361 21345</lparam>
<lparam>Address:5362 21346</lparam>
<lparam>Address:5363 21347</lparam>
<lparam>Address:5364 21348</lparam>
<lparam>Address:5365 21349</lparam>
<lparam>Address:5366 21350</lparam>
<lparam>Address:5367 21351</lparam>
<lparam>Address:5368 21352</lparam>
<lparam>Address:5369 21353</lparam>
<lparam>Address:5370 21360</lparam>
<lparam>Address:5371 21361</lparam>
<lparam>Address:5372 21362</lparam>
<lparam>Address:5373 21363</lparam>
<lparam>Address:5374 21364</lparam>
<lparam>Address:5375 21365</lparam>
<lparam>Address:5376 21366</lparam>
<lparam>Address:5377 21367</lparam>
<lparam>Address:5378 21368</lparam>
<lparam>Address:5379 21369</lparam>
<lparam>Address:5380 21376</lparam>
<lparam>Address:5381 21377</lparam>
<lparam>Address:5382 21378</lparam>
<lparam>Address:5383 21379</lparam>
<lparam>Address:5384 21380</lparam>
<lparam>Address:5385 21381</lparam>
<lparam>Address:5386 21382</lparam>
<lparam>Address:5387 21383</lparam>
<lparam>Address:5388 21384</lparam>
<lparam>Address:5389 21385</lparam>
<lparam>Address:5390 21392</lparam>
<lparam>Address:5391 21393</lparam>
<lparam>Address:5392 21394</lparam>
<lparam>Address:5393 21395</lparam>
<lparam>Address:5394 21396</lparam>
<lparam>Address:5395 21397</lparam>
<lparam>Address:5396 21398</lparam>
<lparam>Address:5397 21399</lparam>
<lparam>Address:5398 21400</lparam>
<lparam>Address:5399 21401</lparam>
<lparam>Address:5400 21504</lparam>
<lparam>Address:5401 21505</lparam>
<lparam>Address:5402 21506</lparam>
<lparam>Address:5403 21507</lparam>
<lparam>Address:5404 21508</lparam>
<lparam>Address:5405 21509</lparam>
<lparam>Address:5406 21510</lparam>
<lparam>Address:5407 21511</lparam>
<lparam>Address:5408 21512</lparam>
<lparam>Address:5409 21513</lparam>
<lparam>Address:5410 21520</lparam>
<lparam>Address:5411 21521</lparam>
<lparam>Address:5412 21522</lparam>
<lparam>Address:5413 21523</lparam>
<lparam>Address:5414 21524</lparam>
<lparam>Address:5415 21525</lparam>
<lparam>Address:5416 21526</lparam>
<lparam>Address:5417 21527</lparam>
<lparam>Address:5418 21528</lparam>
<lparam>Address:5419 21529</lparam>
<lparam>Address:5420 21536</lparam>
<lparam>Address:5421 21537</lparam>
<lparam>Address:5422 21538</lparam>
<lparam>Address:5423 21539</lparam>
<lparam>Address:5424 21540</lparam>
<lparam>Address:5425 21541</lparam>
<lparam>Address:5426 21542</lparam>
<lparam>Address:5427 21543</lparam>
<lparam>Address:5428 21544</lparam>
<lparam>Address:5429 21545</lparam>
<lparam>Address:5430 21552</lparam>
<lparam>Address:5431 21553</lparam>
<lparam>Address:5432 21554</lparam>
<lparam>Address:5433 21555</lparam>
<lparam>Address:5434 21556</lparam>
<lparam>Address:5435 21557</lparam>
<lparam>Address:5436 21558</lparam>
<lparam>Address:5437 21559</lparam>
<lparam>Address:5438 21560</lparam>
<lparam>Address:5439 21561</lparam>
<lparam>Address:5440 21568</lparam>
<lparam>Address:5441 21569</lparam>
<lparam>Address:5442 21570</lparam>
<lparam>Address:5443 21571</lparam>
<lparam>Address:5444 21572</lparam>
<lparam>Address:5445 21573</lparam>
<lparam>Address:5446 21574</lparam>
<lparam>Address:5447 21575</lparam>
<lparam>Address:5448 21576</lparam>
<lparam>Address:5449 21577</lparam>
<lparam>Address:5450 21584</lparam>
<lparam>Address:5451 21585</lparam>
<lparam>Address:5452 21586</lparam>
<lparam>Address:5453 21587</lparam>
<lparam>Address:5454 21588</lparam>
<lparam>Address:5455 21589</lparam>
<lparam>Address:5456 21590</lparam>
<lparam>Address:5457 21591</lparam>
<lparam>Address:5458 21592</lparam>
<lparam>Address:5459 21593</lparam>
<lparam>Address:5460 21600</lparam>
<lparam>Address:5461 21601</lparam>
<lparam>Address:5462 21602</lparam>
<lparam>Address:5463 21603</lparam>
<lparam>Address:5464 21604</lparam>
<lparam>Address:5465 21605</lparam>
<lparam>Address:5466 21606</lparam>
<lparam>Address:5467 21607</lparam>
<lparam>Address:5468 21608</lparam>
<lparam>Address:5469 21609</lparam>
<lparam>Address:5470 21616</lparam>
<lparam>Address:5471 21617</lparam>
<lparam>Address:5472 21618</lparam>
<lparam>Address:5473 21619</lparam>
<lparam>Address:5474 21620</lparam>
<lparam>Address:5475 21621</lparam>
<lparam>Address:5476 21622</lparam>
<lparam>Address:5477 21623</lparam>
<lparam>Address:5478 21624</lparam>
<lparam>Address:5479 21625</lparam>
<lparam>Address:5480 21632</lparam>
<lparam>Address:5481 21633</lparam>
<lparam>Address:5482 21634</lparam>
<lparam>Address:5483 21635</lparam>
<lparam>Address:5484 21636</lparam>
<lparam>Address:5485 21637</lparam>
<lparam>Address:5486 21638</lparam>
<lparam>Address:5487 21639</lparam>
<lparam>Address:5488 21640</lparam>
<lparam>Address:5489 21641</lparam>
<lparam>Address:5490 21648</lparam>
<lparam>Address:5491 21649</lparam>
<lparam>Address:5492 21650</lparam>
<lparam>Address:5493 21651</lparam>
<lparam>Address:5494 21652</lparam>
<lparam>Address:5495 21653</lparam>
<lparam>Address:5496 21654</lparam>
<lparam>Address:5497 21655</lparam>
<lparam>Address:5498 21656</lparam>
<lparam>Address:5499 21657</lparam>
<lparam>Address:5500 21760</lparam>
<lparam>Address:5501 21761</lparam>
<lparam>Address:5502 21762</lparam>
<lparam>Address:5503 21763</lparam>
<lparam>Address:5504 21764</lparam>
<lparam>Address:5505 21765</lparam>
<lparam>Address:5506 21766</lparam>
<lparam>Address:5507 21767</lparam>
<lparam>Address:5508 21768</lparam>
<lparam>Address:5509 21769</lparam>
<lparam>Address:5510 21776</lparam>
<lparam>Address:5511 21777</lparam>
<lparam>Address:5512 21778</lparam>
<lparam>Address:5513 21779</lparam>
<lparam>Address:5514 21780</lparam>
<lparam>Address:5515 21781</lparam>
<lparam>Address:5516 21782</lparam>
<lparam>Address:5517 21783</lparam>
<lparam>Address:5518 21784</lparam>
<lparam>Address:5519 21785</lparam>
<lparam>Address:5520 21792</lparam>
<lparam>Address:5521 21793</lparam>
<lparam>Address:5522 21794</lparam>
<lparam>Address:5523 21795</lparam>
<lparam>Address:5524 21796</lparam>
<lparam>Address:5525 21797</lparam>
<lparam>Address:5526 21798</lparam>
<lparam>Address:5527 21799</lparam>
<lparam>Address:5528 21800</lparam>
<lparam>Address:5529 21801</lparam>
<lparam>Address:5530 21808</lparam>
<lparam>Address:5531 21809</lparam>
<lparam>Address:5532 21810</lparam>
<lparam>Address:5533 21811</lparam>
<lparam>Address:5534 21812</lparam>
<lparam>Address:5535 21813</lparam>
<lparam>Address:5536 21814</lparam>
<lparam>Address:5537 21815</lparam>
<lparam>Address:5538 21816</lparam>
<lparam>Address:5539 21817</lparam>
<lparam>Address:5540 21824</lparam>
<lparam>Address:5541 21825</lparam>
<lparam>Address:5542 21826</lparam>
<lparam>Address:5543 21827</lparam>
<lparam>Address:5544 21828</lparam>
<lparam>Address:5545 21829</lparam>
<lparam>Address:5546 21830</lparam>
<lparam>Address:5547 21831</lparam>
<lparam>Address:5548 21832</lparam>
<lparam>Address:5549 21833</lparam>
<lparam>Address:5550 21840</lparam>
<lparam>Address:5551 21841</lparam>
<lparam>Address:5552 21842</lparam>
<lparam>Address:5553 21843</lparam>
<lparam>Address:5554 21844</lparam>
<lparam>Address:5555 21845</lparam>
<lparam>Address:5556 21846</lparam>
<lparam>Address:5557 21847</lparam>
<lparam>Address:5558 21848</lparam>
<lparam>Address:5559 21849</lparam>
<lparam>Address:5560 21856</lparam>
<lparam>Address:5561 21857</lparam>
<lparam>Address:5562 21858</lparam>
<lparam>Address:5563 21859</lparam>
<lparam>Address:5564 21860</lparam>
<lparam>Address:5565 21861</lparam>
<lparam>Address:5566 21862</lparam>
<lparam>Address:5567 21863</lparam>
<lparam>Address:5568 21864</lparam>
<lparam>Address:5569 21865</lparam>
<lparam>Address:5570 21872</lparam>
<lparam>Address:5571 21873</lparam>
<lparam>Address:5572 21874</lparam>
<lparam>Address:5573 21875</lparam>
<lparam>Address:5574 21876</lparam>
<lparam>Address:5575 21877</lparam>
<lparam>Address:5576 21878</lparam>
<lparam>Address:5577 21879</lparam>
<lparam>Address:5578 21880</lparam>
<lparam>Address:5579 21881</lparam>
<lparam>Address:5580 21888</lparam>
<lparam>Address:5581 21889</lparam>
<lparam>Address:5582 21890</lparam>
<lparam>Address:5583 21891</lparam>
<lparam>Address:5584 21892</lparam>
<lparam>Address:5585 21893</lparam>
<lparam>Address:5586 21894</lparam>
<lparam>Address:5587 21895</lparam>
<lparam>Address:5588 21896</lparam>
<lparam>Address:5589 21897</lparam>
<lparam>Address:5590 21904</lparam>
<lparam>Address:5591 21905</lparam>
<lparam>Address:5592 21906</lparam>
<lparam>Address:5593 21907</lparam>
<lparam>Address:5594 21908</lparam>
<lparam>Address:5595 21909</lparam>
<lparam>Address:5596 21910</lparam>
<lparam>Address:5597 21911</lparam>
<lparam>Address:5598 21912</lparam>
<lparam>Address:5599 21913</lparam>
<lparam>Address:5600 22016</lparam>
<lparam>Address:5601 22017</lparam>
<lparam>Address:5602 22018</lparam>
<lparam>Address:5603 22019</lparam>
<lparam>Address:5604 22020</lparam>
<lparam>Address:5605 22021</lparam>
<lparam>Address:5606 22022</lparam>
<lparam>Address:5607 22023</lparam>
<lparam>Address:5608 22024</lparam>
<lparam>Address:5609 22025</lparam>
<lparam>Address:5610 22032</lparam>
<lparam>Address:5611 22033</lparam>
<lparam>Address:5612 22034</lparam>
<lparam>Address:5613 22035</lparam>
<lparam>Address:5614 22036</lparam>
<lparam>Address:5615 22037</lparam>
<lparam>Address:5616 22038</lparam>
<lparam>Address:5617 22039</lparam>
<lparam>Address:5618 22040</lparam>
<lparam>Address:5619 22041</lparam>
<lparam>Address:5620 22048</lparam>
<lparam>Address:5621 22049</lparam>
<lparam>Address:5622 22050</lparam>
<lparam>Address:5623 22051</lparam>
<lparam>Address:5624 22052</lparam>
<lparam>Address:5625 22053</lparam>
<lparam>Address:5626 22054</lparam>
<lparam>Address:5627 22055</lparam>
<lparam>Address:5628 22056</lparam>
<lparam>Address:5629 22057</lparam>
<lparam>Address:5630 22064</lparam>
<lparam>Address:5631 22065</lparam>
<lparam>Address:5632 22066</lparam>
<lparam>Address:5633 22067</lparam>
<lparam>Address:5634 22068</lparam>
<lparam>Address:5635 22069</lparam>
<lparam>Address:5636 22070</lparam>
<lparam>Address:5637 22071</lparam>
<lparam>Address:5638 22072</lparam>
<lparam>Address:5639 22073</lparam>
<lparam>Address:5640 22080</lparam>
<lparam>Address:5641 22081</lparam>
<lparam>Address:5642 22082</lparam>
<lparam>Address:5643 22083</lparam>
<lparam>Address:5644 22084</lparam>
<lparam>Address:5645 22085</lparam>
<lparam>Address:5646 22086</lparam>
<lparam>Address:5647 22087</lparam>
<lparam>Address:5648 22088</lparam>
<lparam>Address:5649 22089</lparam>
<lparam>Address:5650 22096</lparam>
<lparam>Address:5651 22097</lparam>
<lparam>Address:5652 22098</lparam>
<lparam>Address:5653 22099</lparam>
<lparam>Address:5654 22100</lparam>
<lparam>Address:5655 22101</lparam>
<lparam>Address:5656 22102</lparam>
<lparam>Address:5657 22103</lparam>
<lparam>Address:5658 22104</lparam>
<lparam>Address:5659 22105</lparam>
<lparam>Address:5660 22112</lparam>
<lparam>Address:5661 22113</lparam>
<lparam>Address:5662 22114</lparam>
<lparam>Address:5663 22115</lparam>
<lparam>Address:5664 22116</lparam>
<lparam>Address:5665 22117</lparam>
<lparam>Address:5666 22118</lparam>
<lparam>Address:5667 22119</lparam>
<lparam>Address:5668 22120</lparam>
<lparam>Address:5669 22121</lparam>
<lparam>Address:5670 22128</lparam>
<lparam>Address:5671 22129</lparam>
<lparam>Address:5672 22130</lparam>
<lparam>Address:5673 22131</lparam>
<lparam>Address:5674 22132</lparam>
<lparam>Address:5675 22133</lparam>
<lparam>Address:5676 22134</lparam>
<lparam>Address:5677 22135</lparam>
<lparam>Address:5678 22136</lparam>
<lparam>Address:5679 22137</lparam>
<lparam>Address:5680 22144</lparam>
<lparam>Address:5681 22145</lparam>
<lparam>Address:5682 22146</lparam>
<lparam>Address:5683 22147</lparam>
<lparam>Address:5684 22148</lparam>
<lparam>Address:5685 22149</lparam>
<lparam>Address:5686 22150</lparam>
<lparam>Address:5687 22151</lparam>
<lparam>Address:5688 22152</lparam>
<lparam>Address:5689 22153</lparam>
<lparam>Address:5690 22160</lparam>
<lparam>Address:5691 22161</lparam>
<lparam>Address:5692 22162</lparam>
<lparam>Address:5693 22163</lparam>
<lparam>Address:5694 22164</lparam>
<lparam>Address:5695 22165</lparam>
<lparam>Address:5696 22166</lparam>
<lparam>Address:5697 22167</lparam>
<lparam>Address:5698 22168</lparam>
<lparam>Address:5699 22169</lparam>
<lparam>Address:5700 22272</lparam>
<lparam>Address:5701 22273</lparam>
<lparam>Address:5702 22274</lparam>
<lparam>Address:5703 22275</lparam>
<lparam>Address:5704 22276</lparam>
<lparam>Address:5705 22277</lparam>
<lparam>Address:5706 22278</lparam>
<lparam>Address:5707 22279</lparam>
<lparam>Address:5708 22280</lparam>
<lparam>Address:5709 22281</lparam>
<lparam>Address:5710 22288</lparam>
<lparam>Address:5711 22289</lparam>
<lparam>Address:5712 22290</lparam>
<lparam>Address:5713 22291</lparam>
<lparam>Address:5714 22292</lparam>
<lparam>Address:5715 22293</lparam>
<lparam>Address:5716 22294</lparam>
<lparam>Address:5717 22295</lparam>
<lparam>Address:5718 22296</lparam>
<lparam>Address:5719 22297</lparam>
<lparam>Address:5720 22304</lparam>
<lparam>Address:5721 22305</lparam>
<lparam>Address:5722 22306</lparam>
<lparam>Address:5723 22307</lparam>
<lparam>Address:5724 22308</lparam>
<lparam>Address:5725 22309</lparam>
<lparam>Address:5726 22310</lparam>
<lparam>Address:5727 22311</lparam>
<lparam>Address:5728 22312</lparam>
<lparam>Address:5729 22313</lparam>
<lparam>Address:5730 22320</lparam>
<lparam>Address:5731 22321</lparam>
<lparam>Address:5732 22322</lparam>
<lparam>Address:5733 22323</lparam>
<lparam>Address:5734 22324</lparam>
<lparam>Address:5735 22325</lparam>
<lparam>Address:5736 22326</lparam>
<lparam>Address:5737 22327</lparam>
<lparam>Address:5738 22328</lparam>
<lparam>Address:5739 22329</lparam>
<lparam>Address:5740 22336</lparam>
<lparam>Address:5741 22337</lparam>
<lparam>Address:5742 22338</lparam>
<lparam>Address:5743 22339</lparam>
<lparam>Address:5744 22340</lparam>
<lparam>Address:5745 22341</lparam>
<lparam>Address:5746 22342</lparam>
<lparam>Address:5747 22343</lparam>
<lparam>Address:5748 22344</lparam>
<lparam>Address:5749 22345</lparam>
<lparam>Address:5750 22352</lparam>
<lparam>Address:5751 22353</lparam>
<lparam>Address:5752 22354</lparam>
<lparam>Address:5753 22355</lparam>
<lparam>Address:5754 22356</lparam>
<lparam>Address:5755 22357</lparam>
<lparam>Address:5756 22358</lparam>
<lparam>Address:5757 22359</lparam>
<lparam>Address:5758 22360</lparam>
<lparam>Address:5759 22361</lparam>
<lparam>Address:5760 22368</lparam>
<lparam>Address:5761 22369</lparam>
<lparam>Address:5762 22370</lparam>
<lparam>Address:5763 22371</lparam>
<lparam>Address:5764 22372</lparam>
<lparam>Address:5765 22373</lparam>
<lparam>Address:5766 22374</lparam>
<lparam>Address:5767 22375</lparam>
<lparam>Address:5768 22376</lparam>
<lparam>Address:5769 22377</lparam>
<lparam>Address:5770 22384</lparam>
<lparam>Address:5771 22385</lparam>
<lparam>Address:5772 22386</lparam>
<lparam>Address:5773 22387</lparam>
<lparam>Address:5774 22388</lparam>
<lparam>Address:5775 22389</lparam>
<lparam>Address:5776 22390</lparam>
<lparam>Address:5777 22391</lparam>
<lparam>Address:5778 22392</lparam>
<lparam>Address:5779 22393</lparam>
<lparam>Address:5780 22400</lparam>
<lparam>Address:5781 22401</lparam>
<lparam>Address:5782 22402</lparam>
<lparam>Address:5783 22403</lparam>
<lparam>Address:5784 22404</lparam>
<lparam>Address:5785 22405</lparam>
<lparam>Address:5786 22406</lparam>
<lparam>Address:5787 22407</lparam>
<lparam>Address:5788 22408</lparam>
<lparam>Address:5789 22409</lparam>
<lparam>Address:5790 22416</lparam>
<lparam>Address:5791 22417</lparam>
<lparam>Address:5792 22418</lparam>
<lparam>Address:5793 22419</lparam>
<lparam>Address:5794 22420</lparam>
<lparam>Address:5795 22421</lparam>
<lparam>Address:5796 22422</lparam>
<lparam>Address:5797 22423</lparam>
<lparam>Address:5798 22424</lparam>
<lparam>Address:5799 22425</lparam>
<lparam>Address:5800 22528</lparam>
<lparam>Address:5801 22529</lparam>
<lparam>Address:5802 22530</lparam>
<lparam>Address:5803 22531</lparam>
<lparam>Address:5804 22532</lparam>
<lparam>Address:5805 22533</lparam>
<lparam>Address:5806 22534</lparam>
<lparam>Address:5807 22535</lparam>
<lparam>Address:5808 22536</lparam>
<lparam>Address:5809 22537</lparam>
<lparam>Address:5810 22544</lparam>
<lparam>Address:5811 22545</lparam>
<lparam>Address:5812 22546</lparam>
<lparam>Address:5813 22547</lparam>
<lparam>Address:5814 22548</lparam>
<lparam>Address:5815 22549</lparam>
<lparam>Address:5816 22550</lparam>
<lparam>Address:5817 22551</lparam>
<lparam>Address:5818 22552</lparam>
<lparam>Address:5819 22553</lparam>
<lparam>Address:5820 22560</lparam>
<lparam>Address:5821 22561</lparam>
<lparam>Address:5822 22562</lparam>
<lparam>Address:5823 22563</lparam>
<lparam>Address:5824 22564</lparam>
<lparam>Address:5825 22565</lparam>
<lparam>Address:5826 22566</lparam>
<lparam>Address:5827 22567</lparam>
<lparam>Address:5828 22568</lparam>
<lparam>Address:5829 22569</lparam>
<lparam>Address:5830 22576</lparam>
<lparam>Address:5831 22577</lparam>
<lparam>Address:5832 22578</lparam>
<lparam>Address:5833 22579</lparam>
<lparam>Address:5834 22580</lparam>
<lparam>Address:5835 22581</lparam>
<lparam>Address:5836 22582</lparam>
<lparam>Address:5837 22583</lparam>
<lparam>Address:5838 22584</lparam>
<lparam>Address:5839 22585</lparam>
<lparam>Address:5840 22592</lparam>
<lparam>Address:5841 22593</lparam>
<lparam>Address:5842 22594</lparam>
<lparam>Address:5843 22595</lparam>
<lparam>Address:5844 22596</lparam>
<lparam>Address:5845 22597</lparam>
<lparam>Address:5846 22598</lparam>
<lparam>Address:5847 22599</lparam>
<lparam>Address:5848 22600</lparam>
<lparam>Address:5849 22601</lparam>
<lparam>Address:5850 22608</lparam>
<lparam>Address:5851 22609</lparam>
<lparam>Address:5852 22610</lparam>
<lparam>Address:5853 22611</lparam>
<lparam>Address:5854 22612</lparam>
<lparam>Address:5855 22613</lparam>
<lparam>Address:5856 22614</lparam>
<lparam>Address:5857 22615</lparam>
<lparam>Address:5858 22616</lparam>
<lparam>Address:5859 22617</lparam>
<lparam>Address:5860 22624</lparam>
<lparam>Address:5861 22625</lparam>
<lparam>Address:5862 22626</lparam>
<lparam>Address:5863 22627</lparam>
<lparam>Address:5864 22628</lparam>
<lparam>Address:5865 22629</lparam>
<lparam>Address:5866 22630</lparam>
<lparam>Address:5867 22631</lparam>
<lparam>Address:5868 22632</lparam>
<lparam>Address:5869 22633</lparam>
<lparam>Address:5870 22640</lparam>
<lparam>Address:5871 22641</lparam>
<lparam>Address:5872 22642</lparam>
<lparam>Address:5873 22643</lparam>
<lparam>Address:5874 22644</lparam>
<lparam>Address:5875 22645</lparam>
<lparam>Address:5876 22646</lparam>
<lparam>Address:5877 22647</lparam>
<lparam>Address:5878 22648</lparam>
<lparam>Address:5879 22649</lparam>
<lparam>Address:5880 22656</lparam>
<lparam>Address:5881 22657</lparam>
<lparam>Address:5882 22658</lparam>
<lparam>Address:5883 22659</lparam>
<lparam>Address:5884 22660</lparam>
<lparam>Address:5885 22661</lparam>
<lparam>Address:5886 22662</lparam>
<lparam>Address:5887 22663</lparam>
<lparam>Address:5888 22664</lparam>
<lparam>Address:5889 22665</lparam>
<lparam>Address:5890 22672</lparam>
<lparam>Address:5891 22673</lparam>
<lparam>Address:5892 22674</lparam>
<lparam>Address:5893 22675</lparam>
<lparam>Address:5894 22676</lparam>
<lparam>Address:5895 22677</lparam>
<lparam>Address:5896 22678</lparam>
<lparam>Address:5897 22679</lparam>
<lparam>Address:5898 22680</lparam>
<lparam>Address:5899 22681</lparam>
<lparam>Address:5900 22784</lparam>
<lparam>Address:5901 22785</lparam>
<lparam>Address:5902 22786</lparam>
<lparam>Address:5903 22787</lparam>
<lparam>Address:5904 22788</lparam>
<lparam>Address:5905 22789</lparam>
<lparam>Address:5906 22790</lparam>
<lparam>Address:5907 22791</lparam>
<lparam>Address:5908 22792</lparam>
<lparam>Address:5909 22793</lparam>
<lparam>Address:5910 22800</lparam>
<lparam>Address:5911 22801</lparam>
<lparam>Address:5912 22802</lparam>
<lparam>Address:5913 22803</lparam>
<lparam>Address:5914 22804</lparam>
<lparam>Address:5915 22805</lparam>
<lparam>Address:5916 22806</lparam>
<lparam>Address:5917 22807</lparam>
<lparam>Address:5918 22808</lparam>
<lparam>Address:5919 22809</lparam>
<lparam>Address:5920 22816</lparam>
<lparam>Address:5921 22817</lparam>
<lparam>Address:5922 22818</lparam>
<lparam>Address:5923 22819</lparam>
<lparam>Address:5924 22820</lparam>
<lparam>Address:5925 22821</lparam>
<lparam>Address:5926 22822</lparam>
<lparam>Address:5927 22823</lparam>
<lparam>Address:5928 22824</lparam>
<lparam>Address:5929 22825</lparam>
<lparam>Address:5930 22832</lparam>
<lparam>Address:5931 22833</lparam>
<lparam>Address:5932 22834</lparam>
<lparam>Address:5933 22835</lparam>
<lparam>Address:5934 22836</lparam>
<lparam>Address:5935 22837</lparam>
<lparam>Address:5936 22838</lparam>
<lparam>Address:5937 22839</lparam>
<lparam>Address:5938 22840</lparam>
<lparam>Address:5939 22841</lparam>
<lparam>Address:5940 22848</lparam>
<lparam>Address:5941 22849</lparam>
<lparam>Address:5942 22850</lparam>
<lparam>Address:5943 22851</lparam>
<lparam>Address:5944 22852</lparam>
<lparam>Address:5945 22853</lparam>
<lparam>Address:5946 22854</lparam>
<lparam>Address:5947 22855</lparam>
<lparam>Address:5948 22856</lparam>
<lparam>Address:5949 22857</lparam>
<lparam>Address:5950 22864</lparam>
<lparam>Address:5951 22865</lparam>
<lparam>Address:5952 22866</lparam>
<lparam>Address:5953 22867</lparam>
<lparam>Address:5954 22868</lparam>
<lparam>Address:5955 22869</lparam>
<lparam>Address:5956 22870</lparam>
<lparam>Address:5957 22871</lparam>
<lparam>Address:5958 22872</lparam>
<lparam>Address:5959 22873</lparam>
<lparam>Address:5960 22880</lparam>
<lparam>Address:5961 22881</lparam>
<lparam>Address:5962 22882</lparam>
<lparam>Address:5963 22883</lparam>
<lparam>Address:5964 22884</lparam>
<lparam>Address:5965 22885</lparam>
<lparam>Address:5966 22886</lparam>
<lparam>Address:5967 22887</lparam>
<lparam>Address:5968 22888</lparam>
<lparam>Address:5969 22889</lparam>
<lparam>Address:5970 22896</lparam>
<lparam>Address:5971 22897</lparam>
<lparam>Address:5972 22898</lparam>
<lparam>Address:5973 22899</lparam>
<lparam>Address:5974 22900</lparam>
<lparam>Address:5975 22901</lparam>
<lparam>Address:5976 22902</lparam>
<lparam>Address:5977 22903</lparam>
<lparam>Address:5978 22904</lparam>
<lparam>Address:5979 22905</lparam>
<lparam>Address:5980 22912</lparam>
<lparam>Address:5981 22913</lparam>
<lparam>Address:5982 22914</lparam>
<lparam>Address:5983 22915</lparam>
<lparam>Address:5984 22916</lparam>
<lparam>Address:5985 22917</lparam>
<lparam>Address:5986 22918</lparam>
<lparam>Address:5987 22919</lparam>
<lparam>Address:5988 22920</lparam>
<lparam>Address:5989 22921</lparam>
<lparam>Address:5990 22928</lparam>
<lparam>Address:5991 22929</lparam>
<lparam>Address:5992 22930</lparam>
<lparam>Address:5993 22931</lparam>
<lparam>Address:5994 22932</lparam>
<lparam>Address:5995 22933</lparam>
<lparam>Address:5996 22934</lparam>
<lparam>Address:5997 22935</lparam>
<lparam>Address:5998 22936</lparam>
<lparam>Address:5999 22937</lparam>
<lparam>Address:6000 24576</lparam>
<lparam>Address:6001 24577</lparam>
<lparam>Address:6002 24578</lparam>
<lparam>Address:6003 24579</lparam>
<lparam>Address:6004 24580</lparam>
<lparam>Address:6005 24581</lparam>
<lparam>Address:6006 24582</lparam>
<lparam>Address:6007 24583</lparam>
<lparam>Address:6008 24584</lparam>
<lparam>Address:6009 24585</lparam>
<lparam>Address:6010 24592</lparam>
<lparam>Address:6011 24593</lparam>
<lparam>Address:6012 24594</lparam>
<lparam>Address:6013 24595</lparam>
<lparam>Address:6014 24596</lparam>
<lparam>Address:6015 24597</lparam>
<lparam>Address:6016 24598</lparam>
<lparam>Address:6017 24599</lparam>
<lparam>Address:6018 24600</lparam>
<lparam>Address:6019 24601</lparam>
<lparam>Address:6020 24608</lparam>
<lparam>Address:6021 24609</lparam>
<lparam>Address:6022 24610</lparam>
<lparam>Address:6023 24611</lparam>
<lparam>Address:6024 24612</lparam>
<lparam>Address:6025 24613</lparam>
<lparam>Address:6026 24614</lparam>
<lparam>Address:6027 24615</lparam>
<lparam>Address:6028 24616</lparam>
<lparam>Address:6029 24617</lparam>
<lparam>Address:6030 24624</lparam>
<lparam>Address:6031 24625</lparam>
<lparam>Address:6032 24626</lparam>
<lparam>Address:6033 24627</lparam>
<lparam>Address:6034 24628</lparam>
<lparam>Address:6035 24629</lparam>
<lparam>Address:6036 24630</lparam>
<lparam>Address:6037 24631</lparam>
<lparam>Address:6038 24632</lparam>
<lparam>Address:6039 24633</lparam>
<lparam>Address:6040 24640</lparam>
<lparam>Address:6041 24641</lparam>
<lparam>Address:6042 24642</lparam>
<lparam>Address:6043 24643</lparam>
<lparam>Address:6044 24644</lparam>
<lparam>Address:6045 24645</lparam>
<lparam>Address:6046 24646</lparam>
<lparam>Address:6047 24647</lparam>
<lparam>Address:6048 24648</lparam>
<lparam>Address:6049 24649</lparam>
<lparam>Address:6050 24656</lparam>
<lparam>Address:6051 24657</lparam>
<lparam>Address:6052 24658</lparam>
<lparam>Address:6053 24659</lparam>
<lparam>Address:6054 24660</lparam>
<lparam>Address:6055 24661</lparam>
<lparam>Address:6056 24662</lparam>
<lparam>Address:6057 24663</lparam>
<lparam>Address:6058 24664</lparam>
<lparam>Address:6059 24665</lparam>
<lparam>Address:6060 24672</lparam>
<lparam>Address:6061 24673</lparam>
<lparam>Address:6062 24674</lparam>
<lparam>Address:6063 24675</lparam>
<lparam>Address:6064 24676</lparam>
<lparam>Address:6065 24677</lparam>
<lparam>Address:6066 24678</lparam>
<lparam>Address:6067 24679</lparam>
<lparam>Address:6068 24680</lparam>
<lparam>Address:6069 24681</lparam>
<lparam>Address:6070 24688</lparam>
<lparam>Address:6071 24689</lparam>
<lparam>Address:6072 24690</lparam>
<lparam>Address:6073 24691</lparam>
<lparam>Address:6074 24692</lparam>
<lparam>Address:6075 24693</lparam>
<lparam>Address:6076 24694</lparam>
<lparam>Address:6077 24695</lparam>
<lparam>Address:6078 24696</lparam>
<lparam>Address:6079 24697</lparam>
<lparam>Address:6080 24704</lparam>
<lparam>Address:6081 24705</lparam>
<lparam>Address:6082 24706</lparam>
<lparam>Address:6083 24707</lparam>
<lparam>Address:6084 24708</lparam>
<lparam>Address:6085 24709</lparam>
<lparam>Address:6086 24710</lparam>
<lparam>Address:6087 24711</lparam>
<lparam>Address:6088 24712</lparam>
<lparam>Address:6089 24713</lparam>
<lparam>Address:6090 24720</lparam>
<lparam>Address:6091 24721</lparam>
<lparam>Address:6092 24722</lparam>
<lparam>Address:6093 24723</lparam>
<lparam>Address:6094 24724</lparam>
<lparam>Address:6095 24725</lparam>
<lparam>Address:6096 24726</lparam>
<lparam>Address:6097 24727</lparam>
<lparam>Address:6098 24728</lparam>
<lparam>Address:6099 24729</lparam>
<lparam>Address:6100 24832</lparam>
<lparam>Address:6101 24833</lparam>
<lparam>Address:6102 24834</lparam>
<lparam>Address:6103 24835</lparam>
<lparam>Address:6104 24836</lparam>
<lparam>Address:6105 24837</lparam>
<lparam>Address:6106 24838</lparam>
<lparam>Address:6107 24839</lparam>
<lparam>Address:6108 24840</lparam>
<lparam>Address:6109 24841</lparam>
<lparam>Address:6110 24848</lparam>
<lparam>Address:6111 24849</lparam>
<lparam>Address:6112 24850</lparam>
<lparam>Address:6113 24851</lparam>
<lparam>Address:6114 24852</lparam>
<lparam>Address:6115 24853</lparam>
<lparam>Address:6116 24854</lparam>
<lparam>Address:6117 24855</lparam>
<lparam>Address:6118 24856</lparam>
<lparam>Address:6119 24857</lparam>
<lparam>Address:6120 24864</lparam>
<lparam>Address:6121 24865</lparam>
<lparam>Address:6122 24866</lparam>
<lparam>Address:6123 24867</lparam>
<lparam>Address:6124 24868</lparam>
<lparam>Address:6125 24869</lparam>
<lparam>Address:6126 24870</lparam>
<lparam>Address:6127 24871</lparam>
<lparam>Address:6128 24872</lparam>
<lparam>Address:6129 24873</lparam>
<lparam>Address:6130 24880</lparam>
<lparam>Address:6131 24881</lparam>
<lparam>Address:6132 24882</lparam>
<lparam>Address:6133 24883</lparam>
<lparam>Address:6134 24884</lparam>
<lparam>Address:6135 24885</lparam>
<lparam>Address:6136 24886</lparam>
<lparam>Address:6137 24887</lparam>
<lparam>Address:6138 24888</lparam>
<lparam>Address:6139 24889</lparam>
<lparam>Address:6140 24896</lparam>
<lparam>Address:6141 24897</lparam>
<lparam>Address:6142 24898</lparam>
<lparam>Address:6143 24899</lparam>
<lparam>Address:6144 24900</lparam>
<lparam>Address:6145 24901</lparam>
<lparam>Address:6146 24902</lparam>
<lparam>Address:6147 24903</lparam>
<lparam>Address:6148 24904</lparam>
<lparam>Address:6149 24905</lparam>
<lparam>Address:6150 24912</lparam>
<lparam>Address:6151 24913</lparam>
<lparam>Address:6152 24914</lparam>
<lparam>Address:6153 24915</lparam>
<lparam>Address:6154 24916</lparam>
<lparam>Address:6155 24917</lparam>
<lparam>Address:6156 24918</lparam>
<lparam>Address:6157 24919</lparam>
<lparam>Address:6158 24920</lparam>
<lparam>Address:6159 24921</lparam>
<lparam>Address:6160 24928</lparam>
<lparam>Address:6161 24929</lparam>
<lparam>Address:6162 24930</lparam>
<lparam>Address:6163 24931</lparam>
<lparam>Address:6164 24932</lparam>
<lparam>Address:6165 24933</lparam>
<lparam>Address:6166 24934</lparam>
<lparam>Address:6167 24935</lparam>
<lparam>Address:6168 24936</lparam>
<lparam>Address:6169 24937</lparam>
<lparam>Address:6170 24944</lparam>
<lparam>Address:6171 24945</lparam>
<lparam>Address:6172 24946</lparam>
<lparam>Address:6173 24947</lparam>
<lparam>Address:6174 24948</lparam>
<lparam>Address:6175 24949</lparam>
<lparam>Address:6176 24950</lparam>
<lparam>Address:6177 24951</lparam>
<lparam>Address:6178 24952</lparam>
<lparam>Address:6179 24953</lparam>
<lparam>Address:6180 24960</lparam>
<lparam>Address:6181 24961</lparam>
<lparam>Address:6182 24962</lparam>
<lparam>Address:6183 24963</lparam>
<lparam>Address:6184 24964</lparam>
<lparam>Address:6185 24965</lparam>
<lparam>Address:6186 24966</lparam>
<lparam>Address:6187 24967</lparam>
<lparam>Address:6188 24968</lparam>
<lparam>Address:6189 24969</lparam>
<lparam>Address:6190 24976</lparam>
<lparam>Address:6191 24977</lparam>
<lparam>Address:6192 24978</lparam>
<lparam>Address:6193 24979</lparam>
<lparam>Address:6194 24980</lparam>
<lparam>Address:6195 24981</lparam>
<lparam>Address:6196 24982</lparam>
<lparam>Address:6197 24983</lparam>
<lparam>Address:6198 24984</lparam>
<lparam>Address:6199 24985</lparam>
<lparam>Address:6200 25088</lparam>
<lparam>Address:6201 25089</lparam>
<lparam>Address:6202 25090</lparam>
<lparam>Address:6203 25091</lparam>
<lparam>Address:6204 25092</lparam>
<lparam>Address:6205 25093</lparam>
<lparam>Address:6206 25094</lparam>
<lparam>Address:6207 25095</lparam>
<lparam>Address:6208 25096</lparam>
<lparam>Address:6209 25097</lparam>
<lparam>Address:6210 25104</lparam>
<lparam>Address:6211 25105</lparam>
<lparam>Address:6212 25106</lparam>
<lparam>Address:6213 25107</lparam>
<lparam>Address:6214 25108</lparam>
<lparam>Address:6215 25109</lparam>
<lparam>Address:6216 25110</lparam>
<lparam>Address:6217 25111</lparam>
<lparam>Address:6218 25112</lparam>
<lparam>Address:6219 25113</lparam>
<lparam>Address:6220 25120</lparam>
<lparam>Address:6221 25121</lparam>
<lparam>Address:6222 25122</lparam>
<lparam>Address:6223 25123</lparam>
<lparam>Address:6224 25124</lparam>
<lparam>Address:6225 25125</lparam>
<lparam>Address:6226 25126</lparam>
<lparam>Address:6227 25127</lparam>
<lparam>Address:6228 25128</lparam>
<lparam>Address:6229 25129</lparam>
<lparam>Address:6230 25136</lparam>
<lparam>Address:6231 25137</lparam>
<lparam>Address:6232 25138</lparam>
<lparam>Address:6233 25139</lparam>
<lparam>Address:6234 25140</lparam>
<lparam>Address:6235 25141</lparam>
<lparam>Address:6236 25142</lparam>
<lparam>Address:6237 25143</lparam>
<lparam>Address:6238 25144</lparam>
<lparam>Address:6239 25145</lparam>
<lparam>Address:6240 25152</lparam>
<lparam>Address:6241 25153</lparam>
<lparam>Address:6242 25154</lparam>
<lparam>Address:6243 25155</lparam>
<lparam>Address:6244 25156</lparam>
<lparam>Address:6245 25157</lparam>
<lparam>Address:6246 25158</lparam>
<lparam>Address:6247 25159</lparam>
<lparam>Address:6248 25160</lparam>
<lparam>Address:6249 25161</lparam>
<lparam>Address:6250 25168</lparam>
<lparam>Address:6251 25169</lparam>
<lparam>Address:6252 25170</lparam>
<lparam>Address:6253 25171</lparam>
<lparam>Address:6254 25172</lparam>
<lparam>Address:6255 25173</lparam>
<lparam>Address:6256 25174</lparam>
<lparam>Address:6257 25175</lparam>
<lparam>Address:6258 25176</lparam>
<lparam>Address:6259 25177</lparam>
<lparam>Address:6260 25184</lparam>
<lparam>Address:6261 25185</lparam>
<lparam>Address:6262 25186</lparam>
<lparam>Address:6263 25187</lparam>
<lparam>Address:6264 25188</lparam>
<lparam>Address:6265 25189</lparam>
<lparam>Address:6266 25190</lparam>
<lparam>Address:6267 25191</lparam>
<lparam>Address:6268 25192</lparam>
<lparam>Address:6269 25193</lparam>
<lparam>Address:6270 25200</lparam>
<lparam>Address:6271 25201</lparam>
<lparam>Address:6272 25202</lparam>
<lparam>Address:6273 25203</lparam>
<lparam>Address:6274 25204</lparam>
<lparam>Address:6275 25205</lparam>
<lparam>Address:6276 25206</lparam>
<lparam>Address:6277 25207</lparam>
<lparam>Address:6278 25208</lparam>
<lparam>Address:6279 25209</lparam>
<lparam>Address:6280 25216</lparam>
<lparam>Address:6281 25217</lparam>
<lparam>Address:6282 25218</lparam>
<lparam>Address:6283 25219</lparam>
<lparam>Address:6284 25220</lparam>
<lparam>Address:6285 25221</lparam>
<lparam>Address:6286 25222</lparam>
<lparam>Address:6287 25223</lparam>
<lparam>Address:6288 25224</lparam>
<lparam>Address:6289 25225</lparam>
<lparam>Address:6290 25232</lparam>
<lparam>Address:6291 25233</lparam>
<lparam>Address:6292 25234</lparam>
<lparam>Address:6293 25235</lparam>
<lparam>Address:6294 25236</lparam>
<lparam>Address:6295 25237</lparam>
<lparam>Address:6296 25238</lparam>
<lparam>Address:6297 25239</lparam>
<lparam>Address:6298 25240</lparam>
<lparam>Address:6299 25241</lparam>
<lparam>Address:6300 25344</lparam>
<lparam>Address:6301 25345</lparam>
<lparam>Address:6302 25346</lparam>
<lparam>Address:6303 25347</lparam>
<lparam>Address:6304 25348</lparam>
<lparam>Address:6305 25349</lparam>
<lparam>Address:6306 25350</lparam>
<lparam>Address:6307 25351</lparam>
<lparam>Address:6308 25352</lparam>
<lparam>Address:6309 25353</lparam>
<lparam>Address:6310 25360</lparam>
<lparam>Address:6311 25361</lparam>
<lparam>Address:6312 25362</lparam>
<lparam>Address:6313 25363</lparam>
<lparam>Address:6314 25364</lparam>
<lparam>Address:6315 25365</lparam>
<lparam>Address:6316 25366</lparam>
<lparam>Address:6317 25367</lparam>
<lparam>Address:6318 25368</lparam>
<lparam>Address:6319 25369</lparam>
<lparam>Address:6320 25376</lparam>
<lparam>Address:6321 25377</lparam>
<lparam>Address:6322 25378</lparam>
<lparam>Address:6323 25379</lparam>
<lparam>Address:6324 25380</lparam>
<lparam>Address:6325 25381</lparam>
<lparam>Address:6326 25382</lparam>
<lparam>Address:6327 25383</lparam>
<lparam>Address:6328 25384</lparam>
<lparam>Address:6329 25385</lparam>
<lparam>Address:6330 25392</lparam>
<lparam>Address:6331 25393</lparam>
<lparam>Address:6332 25394</lparam>
<lparam>Address:6333 25395</lparam>
<lparam>Address:6334 25396</lparam>
<lparam>Address:6335 25397</lparam>
<lparam>Address:6336 25398</lparam>
<lparam>Address:6337 25399</lparam>
<lparam>Address:6338 25400</lparam>
<lparam>Address:6339 25401</lparam>
<lparam>Address:6340 25408</lparam>
<lparam>Address:6341 25409</lparam>
<lparam>Address:6342 25410</lparam>
<lparam>Address:6343 25411</lparam>
<lparam>Address:6344 25412</lparam>
<lparam>Address:6345 25413</lparam>
<lparam>Address:6346 25414</lparam>
<lparam>Address:6347 25415</lparam>
<lparam>Address:6348 25416</lparam>
<lparam>Address:6349 25417</lparam>
<lparam>Address:6350 25424</lparam>
<lparam>Address:6351 25425</lparam>
<lparam>Address:6352 25426</lparam>
<lparam>Address:6353 25427</lparam>
<lparam>Address:6354 25428</lparam>
<lparam>Address:6355 25429</lparam>
<lparam>Address:6356 25430</lparam>
<lparam>Address:6357 25431</lparam>
<lparam>Address:6358 25432</lparam>
<lparam>Address:6359 25433</lparam>
<lparam>Address:6360 25440</lparam>
<lparam>Address:6361 25441</lparam>
<lparam>Address:6362 25442</lparam>
<lparam>Address:6363 25443</lparam>
<lparam>Address:6364 25444</lparam>
<lparam>Address:6365 25445</lparam>
<lparam>Address:6366 25446</lparam>
<lparam>Address:6367 25447</lparam>
<lparam>Address:6368 25448</lparam>
<lparam>Address:6369 25449</lparam>
<lparam>Address:6370 25456</lparam>
<lparam>Address:6371 25457</lparam>
<lparam>Address:6372 25458</lparam>
<lparam>Address:6373 25459</lparam>
<lparam>Address:6374 25460</lparam>
<lparam>Address:6375 25461</lparam>
<lparam>Address:6376 25462</lparam>
<lparam>Address:6377 25463</lparam>
<lparam>Address:6378 25464</lparam>
<lparam>Address:6379 25465</lparam>
<lparam>Address:6380 25472</lparam>
<lparam>Address:6381 25473</lparam>
<lparam>Address:6382 25474</lparam>
<lparam>Address:6383 25475</lparam>
<lparam>Address:6384 25476</lparam>
<lparam>Address:6385 25477</lparam>
<lparam>Address:6386 25478</lparam>
<lparam>Address:6387 25479</lparam>
<lparam>Address:6388 25480</lparam>
<lparam>Address:6389 25481</lparam>
<lparam>Address:6390 25488</lparam>
<lparam>Address:6391 25489</lparam>
<lparam>Address:6392 25490</lparam>
<lparam>Address:6393 25491</lparam>
<lparam>Address:6394 25492</lparam>
<lparam>Address:6395 25493</lparam>
<lparam>Address:6396 25494</lparam>
<lparam>Address:6397 25495</lparam>
<lparam>Address:6398 25496</lparam>
<lparam>Address:6399 25497</lparam>
<lparam>Address:6400 25600</lparam>
<lparam>Address:6401 25601</lparam>
<lparam>Address:6402 25602</lparam>
<lparam>Address:6403 25603</lparam>
<lparam>Address:6404 25604</lparam>
<lparam>Address:6405 25605</lparam>
<lparam>Address:6406 25606</lparam>
<lparam>Address:6407 25607</lparam>
<lparam>Address:6408 25608</lparam>
<lparam>Address:6409 25609</lparam>
<lparam>Address:6410 25616</lparam>
<lparam>Address:6411 25617</lparam>
<lparam>Address:6412 25618</lparam>
<lparam>Address:6413 25619</lparam>
<lparam>Address:6414 25620</lparam>
<lparam>Address:6415 25621</lparam>
<lparam>Address:6416 25622</lparam>
<lparam>Address:6417 25623</lparam>
<lparam>Address:6418 25624</lparam>
<lparam>Address:6419 25625</lparam>
<lparam>Address:6420 25632</lparam>
<lparam>Address:6421 25633</lparam>
<lparam>Address:6422 25634</lparam>
<lparam>Address:6423 25635</lparam>
<lparam>Address:6424 25636</lparam>
<lparam>Address:6425 25637</lparam>
<lparam>Address:6426 25638</lparam>
<lparam>Address:6427 25639</lparam>
<lparam>Address:6428 25640</lparam>
<lparam>Address:6429 25641</lparam>
<lparam>Address:6430 25648</lparam>
<lparam>Address:6431 25649</lparam>
<lparam>Address:6432 25650</lparam>
<lparam>Address:6433 25651</lparam>
<lparam>Address:6434 25652</lparam>
<lparam>Address:6435 25653</lparam>
<lparam>Address:6436 25654</lparam>
<lparam>Address:6437 25655</lparam>
<lparam>Address:6438 25656</lparam>
<lparam>Address:6439 25657</lparam>
<lparam>Address:6440 25664</lparam>
<lparam>Address:6441 25665</lparam>
<lparam>Address:6442 25666</lparam>
<lparam>Address:6443 25667</lparam>
<lparam>Address:6444 25668</lparam>
<lparam>Address:6445 25669</lparam>
<lparam>Address:6446 25670</lparam>
<lparam>Address:6447 25671</lparam>
<lparam>Address:6448 25672</lparam>
<lparam>Address:6449 25673</lparam>
<lparam>Address:6450 25680</lparam>
<lparam>Address:6451 25681</lparam>
<lparam>Address:6452 25682</lparam>
<lparam>Address:6453 25683</lparam>
<lparam>Address:6454 25684</lparam>
<lparam>Address:6455 25685</lparam>
<lparam>Address:6456 25686</lparam>
<lparam>Address:6457 25687</lparam>
<lparam>Address:6458 25688</lparam>
<lparam>Address:6459 25689</lparam>
<lparam>Address:6460 25696</lparam>
<lparam>Address:6461 25697</lparam>
<lparam>Address:6462 25698</lparam>
<lparam>Address:6463 25699</lparam>
<lparam>Address:6464 25700</lparam>
<lparam>Address:6465 25701</lparam>
<lparam>Address:6466 25702</lparam>
<lparam>Address:6467 25703</lparam>
<lparam>Address:6468 25704</lparam>
<lparam>Address:6469 25705</lparam>
<lparam>Address:6470 25712</lparam>
<lparam>Address:6471 25713</lparam>
<lparam>Address:6472 25714</lparam>
<lparam>Address:6473 25715</lparam>
<lparam>Address:6474 25716</lparam>
<lparam>Address:6475 25717</lparam>
<lparam>Address:6476 25718</lparam>
<lparam>Address:6477 25719</lparam>
<lparam>Address:6478 25720</lparam>
<lparam>Address:6479 25721</lparam>
<lparam>Address:6480 25728</lparam>
<lparam>Address:6481 25729</lparam>
<lparam>Address:6482 25730</lparam>
<lparam>Address:6483 25731</lparam>
<lparam>Address:6484 25732</lparam>
<lparam>Address:6485 25733</lparam>
<lparam>Address:6486 25734</lparam>
<lparam>Address:6487 25735</lparam>
<lparam>Address:6488 25736</lparam>
<lparam>Address:6489 25737</lparam>
<lparam>Address:6490 25744</lparam>
<lparam>Address:6491 25745</lparam>
<lparam>Address:6492 25746</lparam>
<lparam>Address:6493 25747</lparam>
<lparam>Address:6494 25748</lparam>
<lparam>Address:6495 25749</lparam>
<lparam>Address:6496 25750</lparam>
<lparam>Address:6497 25751</lparam>
<lparam>Address:6498 25752</lparam>
<lparam>Address:6499 25753</lparam>
<lparam>Address:6500 25856</lparam>
<lparam>Address:6501 25857</lparam>
<lparam>Address:6502 25858</lparam>
<lparam>Address:6503 25859</lparam>
<lparam>Address:6504 25860</lparam>
<lparam>Address:6505 25861</lparam>
<lparam>Address:6506 25862</lparam>
<lparam>Address:6507 25863</lparam>
<lparam>Address:6508 25864</lparam>
<lparam>Address:6509 25865</lparam>
<lparam>Address:6510 25872</lparam>
<lparam>Address:6511 25873</lparam>
<lparam>Address:6512 25874</lparam>
<lparam>Address:6513 25875</lparam>
<lparam>Address:6514 25876</lparam>
<lparam>Address:6515 25877</lparam>
<lparam>Address:6516 25878</lparam>
<lparam>Address:6517 25879</lparam>
<lparam>Address:6518 25880</lparam>
<lparam>Address:6519 25881</lparam>
<lparam>Address:6520 25888</lparam>
<lparam>Address:6521 25889</lparam>
<lparam>Address:6522 25890</lparam>
<lparam>Address:6523 25891</lparam>
<lparam>Address:6524 25892</lparam>
<lparam>Address:6525 25893</lparam>
<lparam>Address:6526 25894</lparam>
<lparam>Address:6527 25895</lparam>
<lparam>Address:6528 25896</lparam>
<lparam>Address:6529 25897</lparam>
<lparam>Address:6530 25904</lparam>
<lparam>Address:6531 25905</lparam>
<lparam>Address:6532 25906</lparam>
<lparam>Address:6533 25907</lparam>
<lparam>Address:6534 25908</lparam>
<lparam>Address:6535 25909</lparam>
<lparam>Address:6536 25910</lparam>
<lparam>Address:6537 25911</lparam>
<lparam>Address:6538 25912</lparam>
<lparam>Address:6539 25913</lparam>
<lparam>Address:6540 25920</lparam>
<lparam>Address:6541 25921</lparam>
<lparam>Address:6542 25922</lparam>
<lparam>Address:6543 25923</lparam>
<lparam>Address:6544 25924</lparam>
<lparam>Address:6545 25925</lparam>
<lparam>Address:6546 25926</lparam>
<lparam>Address:6547 25927</lparam>
<lparam>Address:6548 25928</lparam>
<lparam>Address:6549 25929</lparam>
<lparam>Address:6550 25936</lparam>
<lparam>Address:6551 25937</lparam>
<lparam>Address:6552 25938</lparam>
<lparam>Address:6553 25939</lparam>
<lparam>Address:6554 25940</lparam>
<lparam>Address:6555 25941</lparam>
<lparam>Address:6556 25942</lparam>
<lparam>Address:6557 25943</lparam>
<lparam>Address:6558 25944</lparam>
<lparam>Address:6559 25945</lparam>
<lparam>Address:6560 25952</lparam>
<lparam>Address:6561 25953</lparam>
<lparam>Address:6562 25954</lparam>
<lparam>Address:6563 25955</lparam>
<lparam>Address:6564 25956</lparam>
<lparam>Address:6565 25957</lparam>
<lparam>Address:6566 25958</lparam>
<lparam>Address:6567 25959</lparam>
<lparam>Address:6568 25960</lparam>
<lparam>Address:6569 25961</lparam>
<lparam>Address:6570 25968</lparam>
<lparam>Address:6571 25969</lparam>
<lparam>Address:6572 25970</lparam>
<lparam>Address:6573 25971</lparam>
<lparam>Address:6574 25972</lparam>
<lparam>Address:6575 25973</lparam>
<lparam>Address:6576 25974</lparam>
<lparam>Address:6577 25975</lparam>
<lparam>Address:6578 25976</lparam>
<lparam>Address:6579 25977</lparam>
<lparam>Address:6580 25984</lparam>
<lparam>Address:6581 25985</lparam>
<lparam>Address:6582 25986</lparam>
<lparam>Address:6583 25987</lparam>
<lparam>Address:6584 25988</lparam>
<lparam>Address:6585 25989</lparam>
<lparam>Address:6586 25990</lparam>
<lparam>Address:6587 25991</lparam>
<lparam>Address:6588 25992</lparam>
<lparam>Address:6589 25993</lparam>
<lparam>Address:6590 26000</lparam>
<lparam>Address:6591 26001</lparam>
<lparam>Address:6592 26002</lparam>
<lparam>Address:6593 26003</lparam>
<lparam>Address:6594 26004</lparam>
<lparam>Address:6595 26005</lparam>
<lparam>Address:6596 26006</lparam>
<lparam>Address:6597 26007</lparam>
<lparam>Address:6598 26008</lparam>
<lparam>Address:6599 26009</lparam>
<lparam>Address:6600 26112</lparam>
<lparam>Address:6601 26113</lparam>
<lparam>Address:6602 26114</lparam>
<lparam>Address:6603 26115</lparam>
<lparam>Address:6604 26116</lparam>
<lparam>Address:6605 26117</lparam>
<lparam>Address:6606 26118</lparam>
<lparam>Address:6607 26119</lparam>
<lparam>Address:6608 26120</lparam>
<lparam>Address:6609 26121</lparam>
<lparam>Address:6610 26128</lparam>
<lparam>Address:6611 26129</lparam>
<lparam>Address:6612 26130</lparam>
<lparam>Address:6613 26131</lparam>
<lparam>Address:6614 26132</lparam>
<lparam>Address:6615 26133</lparam>
<lparam>Address:6616 26134</lparam>
<lparam>Address:6617 26135</lparam>
<lparam>Address:6618 26136</lparam>
<lparam>Address:6619 26137</lparam>
<lparam>Address:6620 26144</lparam>
<lparam>Address:6621 26145</lparam>
<lparam>Address:6622 26146</lparam>
<lparam>Address:6623 26147</lparam>
<lparam>Address:6624 26148</lparam>
<lparam>Address:6625 26149</lparam>
<lparam>Address:6626 26150</lparam>
<lparam>Address:6627 26151</lparam>
<lparam>Address:6628 26152</lparam>
<lparam>Address:6629 26153</lparam>
<lparam>Address:6630 26160</lparam>
<lparam>Address:6631 26161</lparam>
<lparam>Address:6632 26162</lparam>
<lparam>Address:6633 26163</lparam>
<lparam>Address:6634 26164</lparam>
<lparam>Address:6635 26165</lparam>
<lparam>Address:6636 26166</lparam>
<lparam>Address:6637 26167</lparam>
<lparam>Address:6638 26168</lparam>
<lparam>Address:6639 26169</lparam>
<lparam>Address:6640 26176</lparam>
<lparam>Address:6641 26177</lparam>
<lparam>Address:6642 26178</lparam>
<lparam>Address:6643 26179</lparam>
<lparam>Address:6644 26180</lparam>
<lparam>Address:6645 26181</lparam>
<lparam>Address:6646 26182</lparam>
<lparam>Address:6647 26183</lparam>
<lparam>Address:6648 26184</lparam>
<lparam>Address:6649 26185</lparam>
<lparam>Address:6650 26192</lparam>
<lparam>Address:6651 26193</lparam>
<lparam>Address:6652 26194</lparam>
<lparam>Address:6653 26195</lparam>
<lparam>Address:6654 26196</lparam>
<lparam>Address:6655 26197</lparam>
<lparam>Address:6656 26198</lparam>
<lparam>Address:6657 26199</lparam>
<lparam>Address:6658 26200</lparam>
<lparam>Address:6659 26201</lparam>
<lparam>Address:6660 26208</lparam>
<lparam>Address:6661 26209</lparam>
<lparam>Address:6662 26210</lparam>
<lparam>Address:6663 26211</lparam>
<lparam>Address:6664 26212</lparam>
<lparam>Address:6665 26213</lparam>
<lparam>Address:6666 26214</lparam>
<lparam>Address:6667 26215</lparam>
<lparam>Address:6668 26216</lparam>
<lparam>Address:6669 26217</lparam>
<lparam>Address:6670 26224</lparam>
<lparam>Address:6671 26225</lparam>
<lparam>Address:6672 26226</lparam>
<lparam>Address:6673 26227</lparam>
<lparam>Address:6674 26228</lparam>
<lparam>Address:6675 26229</lparam>
<lparam>Address:6676 26230</lparam>
<lparam>Address:6677 26231</lparam>
<lparam>Address:6678 26232</lparam>
<lparam>Address:6679 26233</lparam>
<lparam>Address:6680 26240</lparam>
<lparam>Address:6681 26241</lparam>
<lparam>Address:6682 26242</lparam>
<lparam>Address:6683 26243</lparam>
<lparam>Address:6684 26244</lparam>
<lparam>Address:6685 26245</lparam>
<lparam>Address:6686 26246</lparam>
<lparam>Address:6687 26247</lparam>
<lparam>Address:6688 26248</lparam>
<lparam>Address:6689 26249</lparam>
<lparam>Address:6690 26256</lparam>
<lparam>Address:6691 26257</lparam>
<lparam>Address:6692 26258</lparam>
<lparam>Address:6693 26259</lparam>
<lparam>Address:6694 26260</lparam>
<lparam>Address:6695 26261</lparam>
<lparam>Address:6696 26262</lparam>
<lparam>Address:6697 26263</lparam>
<lparam>Address:6698 26264</lparam>
<lparam>Address:6699 26265</lparam>
<lparam>Address:6700 26368</lparam>
<lparam>Address:6701 26369</lparam>
<lparam>Address:6702 26370</lparam>
<lparam>Address:6703 26371</lparam>
<lparam>Address:6704 26372</lparam>
<lparam>Address:6705 26373</lparam>
<lparam>Address:6706 26374</lparam>
<lparam>Address:6707 26375</lparam>
<lparam>Address:6708 26376</lparam>
<lparam>Address:6709 26377</lparam>
<lparam>Address:6710 26384</lparam>
<lparam>Address:6711 26385</lparam>
<lparam>Address:6712 26386</lparam>
<lparam>Address:6713 26387</lparam>
<lparam>Address:6714 26388</lparam>
<lparam>Address:6715 26389</lparam>
<lparam>Address:6716 26390</lparam>
<lparam>Address:6717 26391</lparam>
<lparam>Address:6718 26392</lparam>
<lparam>Address:6719 26393</lparam>
<lparam>Address:6720 26400</lparam>
<lparam>Address:6721 26401</lparam>
<lparam>Address:6722 26402</lparam>
<lparam>Address:6723 26403</lparam>
<lparam>Address:6724 26404</lparam>
<lparam>Address:6725 26405</lparam>
<lparam>Address:6726 26406</lparam>
<lparam>Address:6727 26407</lparam>
<lparam>Address:6728 26408</lparam>
<lparam>Address:6729 26409</lparam>
<lparam>Address:6730 26416</lparam>
<lparam>Address:6731 26417</lparam>
<lparam>Address:6732 26418</lparam>
<lparam>Address:6733 26419</lparam>
<lparam>Address:6734 26420</lparam>
<lparam>Address:6735 26421</lparam>
<lparam>Address:6736 26422</lparam>
<lparam>Address:6737 26423</lparam>
<lparam>Address:6738 26424</lparam>
<lparam>Address:6739 26425</lparam>
<lparam>Address:6740 26432</lparam>
<lparam>Address:6741 26433</lparam>
<lparam>Address:6742 26434</lparam>
<lparam>Address:6743 26435</lparam>
<lparam>Address:6744 26436</lparam>
<lparam>Address:6745 26437</lparam>
<lparam>Address:6746 26438</lparam>
<lparam>Address:6747 26439</lparam>
<lparam>Address:6748 26440</lparam>
<lparam>Address:6749 26441</lparam>
<lparam>Address:6750 26448</lparam>
<lparam>Address:6751 26449</lparam>
<lparam>Address:6752 26450</lparam>
<lparam>Address:6753 26451</lparam>
<lparam>Address:6754 26452</lparam>
<lparam>Address:6755 26453</lparam>
<lparam>Address:6756 26454</lparam>
<lparam>Address:6757 26455</lparam>
<lparam>Address:6758 26456</lparam>
<lparam>Address:6759 26457</lparam>
<lparam>Address:6760 26464</lparam>
<lparam>Address:6761 26465</lparam>
<lparam>Address:6762 26466</lparam>
<lparam>Address:6763 26467</lparam>
<lparam>Address:6764 26468</lparam>
<lparam>Address:6765 26469</lparam>
<lparam>Address:6766 26470</lparam>
<lparam>Address:6767 26471</lparam>
<lparam>Address:6768 26472</lparam>
<lparam>Address:6769 26473</lparam>
<lparam>Address:6770 26480</lparam>
<lparam>Address:6771 26481</lparam>
<lparam>Address:6772 26482</lparam>
<lparam>Address:6773 26483</lparam>
<lparam>Address:6774 26484</lparam>
<lparam>Address:6775 26485</lparam>
<lparam>Address:6776 26486</lparam>
<lparam>Address:6777 26487</lparam>
<lparam>Address:6778 26488</lparam>
<lparam>Address:6779 26489</lparam>
<lparam>Address:6780 26496</lparam>
<lparam>Address:6781 26497</lparam>
<lparam>Address:6782 26498</lparam>
<lparam>Address:6783 26499</lparam>
<lparam>Address:6784 26500</lparam>
<lparam>Address:6785 26501</lparam>
<lparam>Address:6786 26502</lparam>
<lparam>Address:6787 26503</lparam>
<lparam>Address:6788 26504</lparam>
<lparam>Address:6789 26505</lparam>
<lparam>Address:6790 26512</lparam>
<lparam>Address:6791 26513</lparam>
<lparam>Address:6792 26514</lparam>
<lparam>Address:6793 26515</lparam>
<lparam>Address:6794 26516</lparam>
<lparam>Address:6795 26517</lparam>
<lparam>Address:6796 26518</lparam>
<lparam>Address:6797 26519</lparam>
<lparam>Address:6798 26520</lparam>
<lparam>Address:6799 26521</lparam>
<lparam>Address:6800 26624</lparam>
<lparam>Address:6801 26625</lparam>
<lparam>Address:6802 26626</lparam>
<lparam>Address:6803 26627</lparam>
<lparam>Address:6804 26628</lparam>
<lparam>Address:6805 26629</lparam>
<lparam>Address:6806 26630</lparam>
<lparam>Address:6807 26631</lparam>
<lparam>Address:6808 26632</lparam>
<lparam>Address:6809 26633</lparam>
<lparam>Address:6810 26640</lparam>
<lparam>Address:6811 26641</lparam>
<lparam>Address:6812 26642</lparam>
<lparam>Address:6813 26643</lparam>
<lparam>Address:6814 26644</lparam>
<lparam>Address:6815 26645</lparam>
<lparam>Address:6816 26646</lparam>
<lparam>Address:6817 26647</lparam>
<lparam>Address:6818 26648</lparam>
<lparam>Address:6819 26649</lparam>
<lparam>Address:6820 26656</lparam>
<lparam>Address:6821 26657</lparam>
<lparam>Address:6822 26658</lparam>
<lparam>Address:6823 26659</lparam>
<lparam>Address:6824 26660</lparam>
<lparam>Address:6825 26661</lparam>
<lparam>Address:6826 26662</lparam>
<lparam>Address:6827 26663</lparam>
<lparam>Address:6828 26664</lparam>
<lparam>Address:6829 26665</lparam>
<lparam>Address:6830 26672</lparam>
<lparam>Address:6831 26673</lparam>
<lparam>Address:6832 26674</lparam>
<lparam>Address:6833 26675</lparam>
<lparam>Address:6834 26676</lparam>
<lparam>Address:6835 26677</lparam>
<lparam>Address:6836 26678</lparam>
<lparam>Address:6837 26679</lparam>
<lparam>Address:6838 26680</lparam>
<lparam>Address:6839 26681</lparam>
<lparam>Address:6840 26688</lparam>
<lparam>Address:6841 26689</lparam>
<lparam>Address:6842 26690</lparam>
<lparam>Address:6843 26691</lparam>
<lparam>Address:6844 26692</lparam>
<lparam>Address:6845 26693</lparam>
<lparam>Address:6846 26694</lparam>
<lparam>Address:6847 26695</lparam>
<lparam>Address:6848 26696</lparam>
<lparam>Address:6849 26697</lparam>
<lparam>Address:6850 26704</lparam>
<lparam>Address:6851 26705</lparam>
<lparam>Address:6852 26706</lparam>
<lparam>Address:6853 26707</lparam>
<lparam>Address:6854 26708</lparam>
<lparam>Address:6855 26709</lparam>
<lparam>Address:6856 26710</lparam>
<lparam>Address:6857 26711</lparam>
<lparam>Address:6858 26712</lparam>
<lparam>Address:6859 26713</lparam>
<lparam>Address:6860 26720</lparam>
<lparam>Address:6861 26721</lparam>
<lparam>Address:6862 26722</lparam>
<lparam>Address:6863 26723</lparam>
<lparam>Address:6864 26724</lparam>
<lparam>Address:6865 26725</lparam>
<lparam>Address:6866 26726</lparam>
<lparam>Address:6867 26727</lparam>
<lparam>Address:6868 26728</lparam>
<lparam>Address:6869 26729</lparam>
<lparam>Address:6870 26736</lparam>
<lparam>Address:6871 26737</lparam>
<lparam>Address:6872 26738</lparam>
<lparam>Address:6873 26739</lparam>
<lparam>Address:6874 26740</lparam>
<lparam>Address:6875 26741</lparam>
<lparam>Address:6876 26742</lparam>
<lparam>Address:6877 26743</lparam>
<lparam>Address:6878 26744</lparam>
<lparam>Address:6879 26745</lparam>
<lparam>Address:6880 26752</lparam>
<lparam>Address:6881 26753</lparam>
<lparam>Address:6882 26754</lparam>
<lparam>Address:6883 26755</lparam>
<lparam>Address:6884 26756</lparam>
<lparam>Address:6885 26757</lparam>
<lparam>Address:6886 26758</lparam>
<lparam>Address:6887 26759</lparam>
<lparam>Address:6888 26760</lparam>
<lparam>Address:6889 26761</lparam>
<lparam>Address:6890 26768</lparam>
<lparam>Address:6891 26769</lparam>
<lparam>Address:6892 26770</lparam>
<lparam>Address:6893 26771</lparam>
<lparam>Address:6894 26772</lparam>
<lparam>Address:6895 26773</lparam>
<lparam>Address:6896 26774</lparam>
<lparam>Address:6897 26775</lparam>
<lparam>Address:6898 26776</lparam>
<lparam>Address:6899 26777</lparam>
<lparam>Address:6900 26880</lparam>
<lparam>Address:6901 26881</lparam>
<lparam>Address:6902 26882</lparam>
<lparam>Address:6903 26883</lparam>
<lparam>Address:6904 26884</lparam>
<lparam>Address:6905 26885</lparam>
<lparam>Address:6906 26886</lparam>
<lparam>Address:6907 26887</lparam>
<lparam>Address:6908 26888</lparam>
<lparam>Address:6909 26889</lparam>
<lparam>Address:6910 26896</lparam>
<lparam>Address:6911 26897</lparam>
<lparam>Address:6912 26898</lparam>
<lparam>Address:6913 26899</lparam>
<lparam>Address:6914 26900</lparam>
<lparam>Address:6915 26901</lparam>
<lparam>Address:6916 26902</lparam>
<lparam>Address:6917 26903</lparam>
<lparam>Address:6918 26904</lparam>
<lparam>Address:6919 26905</lparam>
<lparam>Address:6920 26912</lparam>
<lparam>Address:6921 26913</lparam>
<lparam>Address:6922 26914</lparam>
<lparam>Address:6923 26915</lparam>
<lparam>Address:6924 26916</lparam>
<lparam>Address:6925 26917</lparam>
<lparam>Address:6926 26918</lparam>
<lparam>Address:6927 26919</lparam>
<lparam>Address:6928 26920</lparam>
<lparam>Address:6929 26921</lparam>
<lparam>Address:6930 26928</lparam>
<lparam>Address:6931 26929</lparam>
<lparam>Address:6932 26930</lparam>
<lparam>Address:6933 26931</lparam>
<lparam>Address:6934 26932</lparam>
<lparam>Address:6935 26933</lparam>
<lparam>Address:6936 26934</lparam>
<lparam>Address:6937 26935</lparam>
<lparam>Address:6938 26936</lparam>
<lparam>Address:6939 26937</lparam>
<lparam>Address:6940 26944</lparam>
<lparam>Address:6941 26945</lparam>
<lparam>Address:6942 26946</lparam>
<lparam>Address:6943 26947</lparam>
<lparam>Address:6944 26948</lparam>
<lparam>Address:6945 26949</lparam>
<lparam>Address:6946 26950</lparam>
<lparam>Address:6947 26951</lparam>
<lparam>Address:6948 26952</lparam>
<lparam>Address:6949 26953</lparam>
<lparam>Address:6950 26960</lparam>
<lparam>Address:6951 26961</lparam>
<lparam>Address:6952 26962</lparam>
<lparam>Address:6953 26963</lparam>
<lparam>Address:6954 26964</lparam>
<lparam>Address:6955 26965</lparam>
<lparam>Address:6956 26966</lparam>
<lparam>Address:6957 26967</lparam>
<lparam>Address:6958 26968</lparam>
<lparam>Address:6959 26969</lparam>
<lparam>Address:6960 26976</lparam>
<lparam>Address:6961 26977</lparam>
<lparam>Address:6962 26978</lparam>
<lparam>Address:6963 26979</lparam>
<lparam>Address:6964 26980</lparam>
<lparam>Address:6965 26981</lparam>
<lparam>Address:6966 26982</lparam>
<lparam>Address:6967 26983</lparam>
<lparam>Address:6968 26984</lparam>
<lparam>Address:6969 26985</lparam>
<lparam>Address:6970 26992</lparam>
<lparam>Address:6971 26993</lparam>
<lparam>Address:6972 26994</lparam>
<lparam>Address:6973 26995</lparam>
<lparam>Address:6974 26996</lparam>
<lparam>Address:6975 26997</lparam>
<lparam>Address:6976 26998</lparam>
<lparam>Address:6977 26999</lparam>
<lparam>Address:6978 27000</lparam>
<lparam>Address:6979 27001</lparam>
<lparam>Address:6980 27008</lparam>
<lparam>Address:6981 27009</lparam>
<lparam>Address:6982 27010</lparam>
<lparam>Address:6983 27011</lparam>
<lparam>Address:6984 27012</lparam>
<lparam>Address:6985 27013</lparam>
<lparam>Address:6986 27014</lparam>
<lparam>Address:6987 27015</lparam>
<lparam>Address:6988 27016</lparam>
<lparam>Address:6989 27017</lparam>
<lparam>Address:6990 27024</lparam>
<lparam>Address:6991 27025</lparam>
<lparam>Address:6992 27026</lparam>
<lparam>Address:6993 27027</lparam>
<lparam>Address:6994 27028</lparam>
<lparam>Address:6995 27029</lparam>
<lparam>Address:6996 27030</lparam>
<lparam>Address:6997 27031</lparam>
<lparam>Address:6998 27032</lparam>
<lparam>Address:6999 27033</lparam>
<lparam>Address:7000 28672</lparam>
<lparam>Address:7001 28673</lparam>
<lparam>Address:7002 28674</lparam>
<lparam>Address:7003 28675</lparam>
<lparam>Address:7004 28676</lparam>
<lparam>Address:7005 28677</lparam>
<lparam>Address:7006 28678</lparam>
<lparam>Address:7007 28679</lparam>
<lparam>Address:7008 28680</lparam>
<lparam>Address:7009 28681</lparam>
<lparam>Address:7010 28688</lparam>
<lparam>Address:7011 28689</lparam>
<lparam>Address:7012 28690</lparam>
<lparam>Address:7013 28691</lparam>
<lparam>Address:7014 28692</lparam>
<lparam>Address:7015 28693</lparam>
<lparam>Address:7016 28694</lparam>
<lparam>Address:7017 28695</lparam>
<lparam>Address:7018 28696</lparam>
<lparam>Address:7019 28697</lparam>
<lparam>Address:7020 28704</lparam>
<lparam>Address:7021 28705</lparam>
<lparam>Address:7022 28706</lparam>
<lparam>Address:7023 28707</lparam>
<lparam>Address:7024 28708</lparam>
<lparam>Address:7025 28709</lparam>
<lparam>Address:7026 28710</lparam>
<lparam>Address:7027 28711</lparam>
<lparam>Address:7028 28712</lparam>
<lparam>Address:7029 28713</lparam>
<lparam>Address:7030 28720</lparam>
<lparam>Address:7031 28721</lparam>
<lparam>Address:7032 28722</lparam>
<lparam>Address:7033 28723</lparam>
<lparam>Address:7034 28724</lparam>
<lparam>Address:7035 28725</lparam>
<lparam>Address:7036 28726</lparam>
<lparam>Address:7037 28727</lparam>
<lparam>Address:7038 28728</lparam>
<lparam>Address:7039 28729</lparam>
<lparam>Address:7040 28736</lparam>
<lparam>Address:7041 28737</lparam>
<lparam>Address:7042 28738</lparam>
<lparam>Address:7043 28739</lparam>
<lparam>Address:7044 28740</lparam>
<lparam>Address:7045 28741</lparam>
<lparam>Address:7046 28742</lparam>
<lparam>Address:7047 28743</lparam>
<lparam>Address:7048 28744</lparam>
<lparam>Address:7049 28745</lparam>
<lparam>Address:7050 28752</lparam>
<lparam>Address:7051 28753</lparam>
<lparam>Address:7052 28754</lparam>
<lparam>Address:7053 28755</lparam>
<lparam>Address:7054 28756</lparam>
<lparam>Address:7055 28757</lparam>
<lparam>Address:7056 28758</lparam>
<lparam>Address:7057 28759</lparam>
<lparam>Address:7058 28760</lparam>
<lparam>Address:7059 28761</lparam>
<lparam>Address:7060 28768</lparam>
<lparam>Address:7061 28769</lparam>
<lparam>Address:7062 28770</lparam>
<lparam>Address:7063 28771</lparam>
<lparam>Address:7064 28772</lparam>
<lparam>Address:7065 28773</lparam>
<lparam>Address:7066 28774</lparam>
<lparam>Address:7067 28775</lparam>
<lparam>Address:7068 28776</lparam>
<lparam>Address:7069 28777</lparam>
<lparam>Address:7070 28784</lparam>
<lparam>Address:7071 28785</lparam>
<lparam>Address:7072 28786</lparam>
<lparam>Address:7073 28787</lparam>
<lparam>Address:7074 28788</lparam>
<lparam>Address:7075 28789</lparam>
<lparam>Address:7076 28790</lparam>
<lparam>Address:7077 28791</lparam>
<lparam>Address:7078 28792</lparam>
<lparam>Address:7079 28793</lparam>
<lparam>Address:7080 28800</lparam>
<lparam>Address:7081 28801</lparam>
<lparam>Address:7082 28802</lparam>
<lparam>Address:7083 28803</lparam>
<lparam>Address:7084 28804</lparam>
<lparam>Address:7085 28805</lparam>
<lparam>Address:7086 28806</lparam>
<lparam>Address:7087 28807</lparam>
<lparam>Address:7088 28808</lparam>
<lparam>Address:7089 28809</lparam>
<lparam>Address:7090 28816</lparam>
<lparam>Address:7091 28817</lparam>
<lparam>Address:7092 28818</lparam>
<lparam>Address:7093 28819</lparam>
<lparam>Address:7094 28820</lparam>
<lparam>Address:7095 28821</lparam>
<lparam>Address:7096 28822</lparam>
<lparam>Address:7097 28823</lparam>
<lparam>Address:7098 28824</lparam>
<lparam>Address:7099 28825</lparam>
<lparam>Address:7100 28928</lparam>
<lparam>Address:7101 28929</lparam>
<lparam>Address:7102 28930</lparam>
<lparam>Address:7103 28931</lparam>
<lparam>Address:7104 28932</lparam>
<lparam>Address:7105 28933</lparam>
<lparam>Address:7106 28934</lparam>
<lparam>Address:7107 28935</lparam>
<lparam>Address:7108 28936</lparam>
<lparam>Address:7109 28937</lparam>
<lparam>Address:7110 28944</lparam>
<lparam>Address:7111 28945</lparam>
<lparam>Address:7112 28946</lparam>
<lparam>Address:7113 28947</lparam>
<lparam>Address:7114 28948</lparam>
<lparam>Address:7115 28949</lparam>
<lparam>Address:7116 28950</lparam>
<lparam>Address:7117 28951</lparam>
<lparam>Address:7118 28952</lparam>
<lparam>Address:7119 28953</lparam>
<lparam>Address:7120 28960</lparam>
<lparam>Address:7121 28961</lparam>
<lparam>Address:7122 28962</lparam>
<lparam>Address:7123 28963</lparam>
<lparam>Address:7124 28964</lparam>
<lparam>Address:7125 28965</lparam>
<lparam>Address:7126 28966</lparam>
<lparam>Address:7127 28967</lparam>
<lparam>Address:7128 28968</lparam>
<lparam>Address:7129 28969</lparam>
<lparam>Address:7130 28976</lparam>
<lparam>Address:7131 28977</lparam>
<lparam>Address:7132 28978</lparam>
<lparam>Address:7133 28979</lparam>
<lparam>Address:7134 28980</lparam>
<lparam>Address:7135 28981</lparam>
<lparam>Address:7136 28982</lparam>
<lparam>Address:7137 28983</lparam>
<lparam>Address:7138 28984</lparam>
<lparam>Address:7139 28985</lparam>
<lparam>Address:7140 28992</lparam>
<lparam>Address:7141 28993</lparam>
<lparam>Address:7142 28994</lparam>
<lparam>Address:7143 28995</lparam>
<lparam>Address:7144 28996</lparam>
<lparam>Address:7145 28997</lparam>
<lparam>Address:7146 28998</lparam>
<lparam>Address:7147 28999</lparam>
<lparam>Address:7148 29000</lparam>
<lparam>Address:7149 29001</lparam>
<lparam>Address:7150 29008</lparam>
<lparam>Address:7151 29009</lparam>
<lparam>Address:7152 29010</lparam>
<lparam>Address:7153 29011</lparam>
<lparam>Address:7154 29012</lparam>
<lparam>Address:7155 29013</lparam>
<lparam>Address:7156 29014</lparam>
<lparam>Address:7157 29015</lparam>
<lparam>Address:7158 29016</lparam>
<lparam>Address:7159 29017</lparam>
<lparam>Address:7160 29024</lparam>
<lparam>Address:7161 29025</lparam>
<lparam>Address:7162 29026</lparam>
<lparam>Address:7163 29027</lparam>
<lparam>Address:7164 29028</lparam>
<lparam>Address:7165 29029</lparam>
<lparam>Address:7166 29030</lparam>
<lparam>Address:7167 29031</lparam>
<lparam>Address:7168 29032</lparam>
<lparam>Address:7169 29033</lparam>
<lparam>Address:7170 29040</lparam>
<lparam>Address:7171 29041</lparam>
<lparam>Address:7172 29042</lparam>
<lparam>Address:7173 29043</lparam>
<lparam>Address:7174 29044</lparam>
<lparam>Address:7175 29045</lparam>
<lparam>Address:7176 29046</lparam>
<lparam>Address:7177 29047</lparam>
<lparam>Address:7178 29048</lparam>
<lparam>Address:7179 29049</lparam>
<lparam>Address:7180 29056</lparam>
<lparam>Address:7181 29057</lparam>
<lparam>Address:7182 29058</lparam>
<lparam>Address:7183 29059</lparam>
<lparam>Address:7184 29060</lparam>
<lparam>Address:7185 29061</lparam>
<lparam>Address:7186 29062</lparam>
<lparam>Address:7187 29063</lparam>
<lparam>Address:7188 29064</lparam>
<lparam>Address:7189 29065</lparam>
<lparam>Address:7190 29072</lparam>
<lparam>Address:7191 29073</lparam>
<lparam>Address:7192 29074</lparam>
<lparam>Address:7193 29075</lparam>
<lparam>Address:7194 29076</lparam>
<lparam>Address:7195 29077</lparam>
<lparam>Address:7196 29078</lparam>
<lparam>Address:7197 29079</lparam>
<lparam>Address:7198 29080</lparam>
<lparam>Address:7199 29081</lparam>
<lparam>Address:7200 29184</lparam>
<lparam>Address:7201 29185</lparam>
<lparam>Address:7202 29186</lparam>
<lparam>Address:7203 29187</lparam>
<lparam>Address:7204 29188</lparam>
<lparam>Address:7205 29189</lparam>
<lparam>Address:7206 29190</lparam>
<lparam>Address:7207 29191</lparam>
<lparam>Address:7208 29192</lparam>
<lparam>Address:7209 29193</lparam>
<lparam>Address:7210 29200</lparam>
<lparam>Address:7211 29201</lparam>
<lparam>Address:7212 29202</lparam>
<lparam>Address:7213 29203</lparam>
<lparam>Address:7214 29204</lparam>
<lparam>Address:7215 29205</lparam>
<lparam>Address:7216 29206</lparam>
<lparam>Address:7217 29207</lparam>
<lparam>Address:7218 29208</lparam>
<lparam>Address:7219 29209</lparam>
<lparam>Address:7220 29216</lparam>
<lparam>Address:7221 29217</lparam>
<lparam>Address:7222 29218</lparam>
<lparam>Address:7223 29219</lparam>
<lparam>Address:7224 29220</lparam>
<lparam>Address:7225 29221</lparam>
<lparam>Address:7226 29222</lparam>
<lparam>Address:7227 29223</lparam>
<lparam>Address:7228 29224</lparam>
<lparam>Address:7229 29225</lparam>
<lparam>Address:7230 29232</lparam>
<lparam>Address:7231 29233</lparam>
<lparam>Address:7232 29234</lparam>
<lparam>Address:7233 29235</lparam>
<lparam>Address:7234 29236</lparam>
<lparam>Address:7235 29237</lparam>
<lparam>Address:7236 29238</lparam>
<lparam>Address:7237 29239</lparam>
<lparam>Address:7238 29240</lparam>
<lparam>Address:7239 29241</lparam>
<lparam>Address:7240 29248</lparam>
<lparam>Address:7241 29249</lparam>
<lparam>Address:7242 29250</lparam>
<lparam>Address:7243 29251</lparam>
<lparam>Address:7244 29252</lparam>
<lparam>Address:7245 29253</lparam>
<lparam>Address:7246 29254</lparam>
<lparam>Address:7247 29255</lparam>
<lparam>Address:7248 29256</lparam>
<lparam>Address:7249 29257</lparam>
<lparam>Address:7250 29264</lparam>
<lparam>Address:7251 29265</lparam>
<lparam>Address:7252 29266</lparam>
<lparam>Address:7253 29267</lparam>
<lparam>Address:7254 29268</lparam>
<lparam>Address:7255 29269</lparam>
<lparam>Address:7256 29270</lparam>
<lparam>Address:7257 29271</lparam>
<lparam>Address:7258 29272</lparam>
<lparam>Address:7259 29273</lparam>
<lparam>Address:7260 29280</lparam>
<lparam>Address:7261 29281</lparam>
<lparam>Address:7262 29282</lparam>
<lparam>Address:7263 29283</lparam>
<lparam>Address:7264 29284</lparam>
<lparam>Address:7265 29285</lparam>
<lparam>Address:7266 29286</lparam>
<lparam>Address:7267 29287</lparam>
<lparam>Address:7268 29288</lparam>
<lparam>Address:7269 29289</lparam>
<lparam>Address:7270 29296</lparam>
<lparam>Address:7271 29297</lparam>
<lparam>Address:7272 29298</lparam>
<lparam>Address:7273 29299</lparam>
<lparam>Address:7274 29300</lparam>
<lparam>Address:7275 29301</lparam>
<lparam>Address:7276 29302</lparam>
<lparam>Address:7277 29303</lparam>
<lparam>Address:7278 29304</lparam>
<lparam>Address:7279 29305</lparam>
<lparam>Address:7280 29312</lparam>
<lparam>Address:7281 29313</lparam>
<lparam>Address:7282 29314</lparam>
<lparam>Address:7283 29315</lparam>
<lparam>Address:7284 29316</lparam>
<lparam>Address:7285 29317</lparam>
<lparam>Address:7286 29318</lparam>
<lparam>Address:7287 29319</lparam>
<lparam>Address:7288 29320</lparam>
<lparam>Address:7289 29321</lparam>
<lparam>Address:7290 29328</lparam>
<lparam>Address:7291 29329</lparam>
<lparam>Address:7292 29330</lparam>
<lparam>Address:7293 29331</lparam>
<lparam>Address:7294 29332</lparam>
<lparam>Address:7295 29333</lparam>
<lparam>Address:7296 29334</lparam>
<lparam>Address:7297 29335</lparam>
<lparam>Address:7298 29336</lparam>
<lparam>Address:7299 29337</lparam>
<lparam>Address:7300 29440</lparam>
<lparam>Address:7301 29441</lparam>
<lparam>Address:7302 29442</lparam>
<lparam>Address:7303 29443</lparam>
<lparam>Address:7304 29444</lparam>
<lparam>Address:7305 29445</lparam>
<lparam>Address:7306 29446</lparam>
<lparam>Address:7307 29447</lparam>
<lparam>Address:7308 29448</lparam>
<lparam>Address:7309 29449</lparam>
<lparam>Address:7310 29456</lparam>
<lparam>Address:7311 29457</lparam>
<lparam>Address:7312 29458</lparam>
<lparam>Address:7313 29459</lparam>
<lparam>Address:7314 29460</lparam>
<lparam>Address:7315 29461</lparam>
<lparam>Address:7316 29462</lparam>
<lparam>Address:7317 29463</lparam>
<lparam>Address:7318 29464</lparam>
<lparam>Address:7319 29465</lparam>
<lparam>Address:7320 29472</lparam>
<lparam>Address:7321 29473</lparam>
<lparam>Address:7322 29474</lparam>
<lparam>Address:7323 29475</lparam>
<lparam>Address:7324 29476</lparam>
<lparam>Address:7325 29477</lparam>
<lparam>Address:7326 29478</lparam>
<lparam>Address:7327 29479</lparam>
<lparam>Address:7328 29480</lparam>
<lparam>Address:7329 29481</lparam>
<lparam>Address:7330 29488</lparam>
<lparam>Address:7331 29489</lparam>
<lparam>Address:7332 29490</lparam>
<lparam>Address:7333 29491</lparam>
<lparam>Address:7334 29492</lparam>
<lparam>Address:7335 29493</lparam>
<lparam>Address:7336 29494</lparam>
<lparam>Address:7337 29495</lparam>
<lparam>Address:7338 29496</lparam>
<lparam>Address:7339 29497</lparam>
<lparam>Address:7340 29504</lparam>
<lparam>Address:7341 29505</lparam>
<lparam>Address:7342 29506</lparam>
<lparam>Address:7343 29507</lparam>
<lparam>Address:7344 29508</lparam>
<lparam>Address:7345 29509</lparam>
<lparam>Address:7346 29510</lparam>
<lparam>Address:7347 29511</lparam>
<lparam>Address:7348 29512</lparam>
<lparam>Address:7349 29513</lparam>
<lparam>Address:7350 29520</lparam>
<lparam>Address:7351 29521</lparam>
<lparam>Address:7352 29522</lparam>
<lparam>Address:7353 29523</lparam>
<lparam>Address:7354 29524</lparam>
<lparam>Address:7355 29525</lparam>
<lparam>Address:7356 29526</lparam>
<lparam>Address:7357 29527</lparam>
<lparam>Address:7358 29528</lparam>
<lparam>Address:7359 29529</lparam>
<lparam>Address:7360 29536</lparam>
<lparam>Address:7361 29537</lparam>
<lparam>Address:7362 29538</lparam>
<lparam>Address:7363 29539</lparam>
<lparam>Address:7364 29540</lparam>
<lparam>Address:7365 29541</lparam>
<lparam>Address:7366 29542</lparam>
<lparam>Address:7367 29543</lparam>
<lparam>Address:7368 29544</lparam>
<lparam>Address:7369 29545</lparam>
<lparam>Address:7370 29552</lparam>
<lparam>Address:7371 29553</lparam>
<lparam>Address:7372 29554</lparam>
<lparam>Address:7373 29555</lparam>
<lparam>Address:7374 29556</lparam>
<lparam>Address:7375 29557</lparam>
<lparam>Address:7376 29558</lparam>
<lparam>Address:7377 29559</lparam>
<lparam>Address:7378 29560</lparam>
<lparam>Address:7379 29561</lparam>
<lparam>Address:7380 29568</lparam>
<lparam>Address:7381 29569</lparam>
<lparam>Address:7382 29570</lparam>
<lparam>Address:7383 29571</lparam>
<lparam>Address:7384 29572</lparam>
<lparam>Address:7385 29573</lparam>
<lparam>Address:7386 29574</lparam>
<lparam>Address:7387 29575</lparam>
<lparam>Address:7388 29576</lparam>
<lparam>Address:7389 29577</lparam>
<lparam>Address:7390 29584</lparam>
<lparam>Address:7391 29585</lparam>
<lparam>Address:7392 29586</lparam>
<lparam>Address:7393 29587</lparam>
<lparam>Address:7394 29588</lparam>
<lparam>Address:7395 29589</lparam>
<lparam>Address:7396 29590</lparam>
<lparam>Address:7397 29591</lparam>
<lparam>Address:7398 29592</lparam>
<lparam>Address:7399 29593</lparam>
<lparam>Address:7400 29696</lparam>
<lparam>Address:7401 29697</lparam>
<lparam>Address:7402 29698</lparam>
<lparam>Address:7403 29699</lparam>
<lparam>Address:7404 29700</lparam>
<lparam>Address:7405 29701</lparam>
<lparam>Address:7406 29702</lparam>
<lparam>Address:7407 29703</lparam>
<lparam>Address:7408 29704</lparam>
<lparam>Address:7409 29705</lparam>
<lparam>Address:7410 29712</lparam>
<lparam>Address:7411 29713</lparam>
<lparam>Address:7412 29714</lparam>
<lparam>Address:7413 29715</lparam>
<lparam>Address:7414 29716</lparam>
<lparam>Address:7415 29717</lparam>
<lparam>Address:7416 29718</lparam>
<lparam>Address:7417 29719</lparam>
<lparam>Address:7418 29720</lparam>
<lparam>Address:7419 29721</lparam>
<lparam>Address:7420 29728</lparam>
<lparam>Address:7421 29729</lparam>
<lparam>Address:7422 29730</lparam>
<lparam>Address:7423 29731</lparam>
<lparam>Address:7424 29732</lparam>
<lparam>Address:7425 29733</lparam>
<lparam>Address:7426 29734</lparam>
<lparam>Address:7427 29735</lparam>
<lparam>Address:7428 29736</lparam>
<lparam>Address:7429 29737</lparam>
<lparam>Address:7430 29744</lparam>
<lparam>Address:7431 29745</lparam>
<lparam>Address:7432 29746</lparam>
<lparam>Address:7433 29747</lparam>
<lparam>Address:7434 29748</lparam>
<lparam>Address:7435 29749</lparam>
<lparam>Address:7436 29750</lparam>
<lparam>Address:7437 29751</lparam>
<lparam>Address:7438 29752</lparam>
<lparam>Address:7439 29753</lparam>
<lparam>Address:7440 29760</lparam>
<lparam>Address:7441 29761</lparam>
<lparam>Address:7442 29762</lparam>
<lparam>Address:7443 29763</lparam>
<lparam>Address:7444 29764</lparam>
<lparam>Address:7445 29765</lparam>
<lparam>Address:7446 29766</lparam>
<lparam>Address:7447 29767</lparam>
<lparam>Address:7448 29768</lparam>
<lparam>Address:7449 29769</lparam>
<lparam>Address:7450 29776</lparam>
<lparam>Address:7451 29777</lparam>
<lparam>Address:7452 29778</lparam>
<lparam>Address:7453 29779</lparam>
<lparam>Address:7454 29780</lparam>
<lparam>Address:7455 29781</lparam>
<lparam>Address:7456 29782</lparam>
<lparam>Address:7457 29783</lparam>
<lparam>Address:7458 29784</lparam>
<lparam>Address:7459 29785</lparam>
<lparam>Address:7460 29792</lparam>
<lparam>Address:7461 29793</lparam>
<lparam>Address:7462 29794</lparam>
<lparam>Address:7463 29795</lparam>
<lparam>Address:7464 29796</lparam>
<lparam>Address:7465 29797</lparam>
<lparam>Address:7466 29798</lparam>
<lparam>Address:7467 29799</lparam>
<lparam>Address:7468 29800</lparam>
<lparam>Address:7469 29801</lparam>
<lparam>Address:7470 29808</lparam>
<lparam>Address:7471 29809</lparam>
<lparam>Address:7472 29810</lparam>
<lparam>Address:7473 29811</lparam>
<lparam>Address:7474 29812</lparam>
<lparam>Address:7475 29813</lparam>
<lparam>Address:7476 29814</lparam>
<lparam>Address:7477 29815</lparam>
<lparam>Address:7478 29816</lparam>
<lparam>Address:7479 29817</lparam>
<lparam>Address:7480 29824</lparam>
<lparam>Address:7481 29825</lparam>
<lparam>Address:7482 29826</lparam>
<lparam>Address:7483 29827</lparam>
<lparam>Address:7484 29828</lparam>
<lparam>Address:7485 29829</lparam>
<lparam>Address:7486 29830</lparam>
<lparam>Address:7487 29831</lparam>
<lparam>Address:7488 29832</lparam>
<lparam>Address:7489 29833</lparam>
<lparam>Address:7490 29840</lparam>
<lparam>Address:7491 29841</lparam>
<lparam>Address:7492 29842</lparam>
<lparam>Address:7493 29843</lparam>
<lparam>Address:7494 29844</lparam>
<lparam>Address:7495 29845</lparam>
<lparam>Address:7496 29846</lparam>
<lparam>Address:7497 29847</lparam>
<lparam>Address:7498 29848</lparam>
<lparam>Address:7499 29849</lparam>
<lparam>Address:7500 29952</lparam>
<lparam>Address:7501 29953</lparam>
<lparam>Address:7502 29954</lparam>
<lparam>Address:7503 29955</lparam>
<lparam>Address:7504 29956</lparam>
<lparam>Address:7505 29957</lparam>
<lparam>Address:7506 29958</lparam>
<lparam>Address:7507 29959</lparam>
<lparam>Address:7508 29960</lparam>
<lparam>Address:7509 29961</lparam>
<lparam>Address:7510 29968</lparam>
<lparam>Address:7511 29969</lparam>
<lparam>Address:7512 29970</lparam>
<lparam>Address:7513 29971</lparam>
<lparam>Address:7514 29972</lparam>
<lparam>Address:7515 29973</lparam>
<lparam>Address:7516 29974</lparam>
<lparam>Address:7517 29975</lparam>
<lparam>Address:7518 29976</lparam>
<lparam>Address:7519 29977</lparam>
<lparam>Address:7520 29984</lparam>
<lparam>Address:7521 29985</lparam>
<lparam>Address:7522 29986</lparam>
<lparam>Address:7523 29987</lparam>
<lparam>Address:7524 29988</lparam>
<lparam>Address:7525 29989</lparam>
<lparam>Address:7526 29990</lparam>
<lparam>Address:7527 29991</lparam>
<lparam>Address:7528 29992</lparam>
<lparam>Address:7529 29993</lparam>
<lparam>Address:7530 30000</lparam>
<lparam>Address:7531 30001</lparam>
<lparam>Address:7532 30002</lparam>
<lparam>Address:7533 30003</lparam>
<lparam>Address:7534 30004</lparam>
<lparam>Address:7535 30005</lparam>
<lparam>Address:7536 30006</lparam>
<lparam>Address:7537 30007</lparam>
<lparam>Address:7538 30008</lparam>
<lparam>Address:7539 30009</lparam>
<lparam>Address:7540 30016</lparam>
<lparam>Address:7541 30017</lparam>
<lparam>Address:7542 30018</lparam>
<lparam>Address:7543 30019</lparam>
<lparam>Address:7544 30020</lparam>
<lparam>Address:7545 30021</lparam>
<lparam>Address:7546 30022</lparam>
<lparam>Address:7547 30023</lparam>
<lparam>Address:7548 30024</lparam>
<lparam>Address:7549 30025</lparam>
<lparam>Address:7550 30032</lparam>
<lparam>Address:7551 30033</lparam>
<lparam>Address:7552 30034</lparam>
<lparam>Address:7553 30035</lparam>
<lparam>Address:7554 30036</lparam>
<lparam>Address:7555 30037</lparam>
<lparam>Address:7556 30038</lparam>
<lparam>Address:7557 30039</lparam>
<lparam>Address:7558 30040</lparam>
<lparam>Address:7559 30041</lparam>
<lparam>Address:7560 30048</lparam>
<lparam>Address:7561 30049</lparam>
<lparam>Address:7562 30050</lparam>
<lparam>Address:7563 30051</lparam>
<lparam>Address:7564 30052</lparam>
<lparam>Address:7565 30053</lparam>
<lparam>Address:7566 30054</lparam>
<lparam>Address:7567 30055</lparam>
<lparam>Address:7568 30056</lparam>
<lparam>Address:7569 30057</lparam>
<lparam>Address:7570 30064</lparam>
<lparam>Address:7571 30065</lparam>
<lparam>Address:7572 30066</lparam>
<lparam>Address:7573 30067</lparam>
<lparam>Address:7574 30068</lparam>
<lparam>Address:7575 30069</lparam>
<lparam>Address:7576 30070</lparam>
<lparam>Address:7577 30071</lparam>
<lparam>Address:7578 30072</lparam>
<lparam>Address:7579 30073</lparam>
<lparam>Address:7580 30080</lparam>
<lparam>Address:7581 30081</lparam>
<lparam>Address:7582 30082</lparam>
<lparam>Address:7583 30083</lparam>
<lparam>Address:7584 30084</lparam>
<lparam>Address:7585 30085</lparam>
<lparam>Address:7586 30086</lparam>
<lparam>Address:7587 30087</lparam>
<lparam>Address:7588 30088</lparam>
<lparam>Address:7589 30089</lparam>
<lparam>Address:7590 30096</lparam>
<lparam>Address:7591 30097</lparam>
<lparam>Address:7592 30098</lparam>
<lparam>Address:7593 30099</lparam>
<lparam>Address:7594 30100</lparam>
<lparam>Address:7595 30101</lparam>
<lparam>Address:7596 30102</lparam>
<lparam>Address:7597 30103</lparam>
<lparam>Address:7598 30104</lparam>
<lparam>Address:7599 30105</lparam>
<lparam>Address:7600 30208</lparam>
<lparam>Address:7601 30209</lparam>
<lparam>Address:7602 30210</lparam>
<lparam>Address:7603 30211</lparam>
<lparam>Address:7604 30212</lparam>
<lparam>Address:7605 30213</lparam>
<lparam>Address:7606 30214</lparam>
<lparam>Address:7607 30215</lparam>
<lparam>Address:7608 30216</lparam>
<lparam>Address:7609 30217</lparam>
<lparam>Address:7610 30224</lparam>
<lparam>Address:7611 30225</lparam>
<lparam>Address:7612 30226</lparam>
<lparam>Address:7613 30227</lparam>
<lparam>Address:7614 30228</lparam>
<lparam>Address:7615 30229</lparam>
<lparam>Address:7616 30230</lparam>
<lparam>Address:7617 30231</lparam>
<lparam>Address:7618 30232</lparam>
<lparam>Address:7619 30233</lparam>
<lparam>Address:7620 30240</lparam>
<lparam>Address:7621 30241</lparam>
<lparam>Address:7622 30242</lparam>
<lparam>Address:7623 30243</lparam>
<lparam>Address:7624 30244</lparam>
<lparam>Address:7625 30245</lparam>
<lparam>Address:7626 30246</lparam>
<lparam>Address:7627 30247</lparam>
<lparam>Address:7628 30248</lparam>
<lparam>Address:7629 30249</lparam>
<lparam>Address:7630 30256</lparam>
<lparam>Address:7631 30257</lparam>
<lparam>Address:7632 30258</lparam>
<lparam>Address:7633 30259</lparam>
<lparam>Address:7634 30260</lparam>
<lparam>Address:7635 30261</lparam>
<lparam>Address:7636 30262</lparam>
<lparam>Address:7637 30263</lparam>
<lparam>Address:7638 30264</lparam>
<lparam>Address:7639 30265</lparam>
<lparam>Address:7640 30272</lparam>
<lparam>Address:7641 30273</lparam>
<lparam>Address:7642 30274</lparam>
<lparam>Address:7643 30275</lparam>
<lparam>Address:7644 30276</lparam>
<lparam>Address:7645 30277</lparam>
<lparam>Address:7646 30278</lparam>
<lparam>Address:7647 30279</lparam>
<lparam>Address:7648 30280</lparam>
<lparam>Address:7649 30281</lparam>
<lparam>Address:7650 30288</lparam>
<lparam>Address:7651 30289</lparam>
<lparam>Address:7652 30290</lparam>
<lparam>Address:7653 30291</lparam>
<lparam>Address:7654 30292</lparam>
<lparam>Address:7655 30293</lparam>
<lparam>Address:7656 30294</lparam>
<lparam>Address:7657 30295</lparam>
<lparam>Address:7658 30296</lparam>
<lparam>Address:7659 30297</lparam>
<lparam>Address:7660 30304</lparam>
<lparam>Address:7661 30305</lparam>
<lparam>Address:7662 30306</lparam>
<lparam>Address:7663 30307</lparam>
<lparam>Address:7664 30308</lparam>
<lparam>Address:7665 30309</lparam>
<lparam>Address:7666 30310</lparam>
<lparam>Address:7667 30311</lparam>
<lparam>Address:7668 30312</lparam>
<lparam>Address:7669 30313</lparam>
<lparam>Address:7670 30320</lparam>
<lparam>Address:7671 30321</lparam>
<lparam>Address:7672 30322</lparam>
<lparam>Address:7673 30323</lparam>
<lparam>Address:7674 30324</lparam>
<lparam>Address:7675 30325</lparam>
<lparam>Address:7676 30326</lparam>
<lparam>Address:7677 30327</lparam>
<lparam>Address:7678 30328</lparam>
<lparam>Address:7679 30329</lparam>
<lparam>Address:7680 30336</lparam>
<lparam>Address:7681 30337</lparam>
<lparam>Address:7682 30338</lparam>
<lparam>Address:7683 30339</lparam>
<lparam>Address:7684 30340</lparam>
<lparam>Address:7685 30341</lparam>
<lparam>Address:7686 30342</lparam>
<lparam>Address:7687 30343</lparam>
<lparam>Address:7688 30344</lparam>
<lparam>Address:7689 30345</lparam>
<lparam>Address:7690 30352</lparam>
<lparam>Address:7691 30353</lparam>
<lparam>Address:7692 30354</lparam>
<lparam>Address:7693 30355</lparam>
<lparam>Address:7694 30356</lparam>
<lparam>Address:7695 30357</lparam>
<lparam>Address:7696 30358</lparam>
<lparam>Address:7697 30359</lparam>
<lparam>Address:7698 30360</lparam>
<lparam>Address:7699 30361</lparam>
<lparam>Address:7700 30464</lparam>
<lparam>Address:7701 30465</lparam>
<lparam>Address:7702 30466</lparam>
<lparam>Address:7703 30467</lparam>
<lparam>Address:7704 30468</lparam>
<lparam>Address:7705 30469</lparam>
<lparam>Address:7706 30470</lparam>
<lparam>Address:7707 30471</lparam>
<lparam>Address:7708 30472</lparam>
<lparam>Address:7709 30473</lparam>
<lparam>Address:7710 30480</lparam>
<lparam>Address:7711 30481</lparam>
<lparam>Address:7712 30482</lparam>
<lparam>Address:7713 30483</lparam>
<lparam>Address:7714 30484</lparam>
<lparam>Address:7715 30485</lparam>
<lparam>Address:7716 30486</lparam>
<lparam>Address:7717 30487</lparam>
<lparam>Address:7718 30488</lparam>
<lparam>Address:7719 30489</lparam>
<lparam>Address:7720 30496</lparam>
<lparam>Address:7721 30497</lparam>
<lparam>Address:7722 30498</lparam>
<lparam>Address:7723 30499</lparam>
<lparam>Address:7724 30500</lparam>
<lparam>Address:7725 30501</lparam>
<lparam>Address:7726 30502</lparam>
<lparam>Address:7727 30503</lparam>
<lparam>Address:7728 30504</lparam>
<lparam>Address:7729 30505</lparam>
<lparam>Address:7730 30512</lparam>
<lparam>Address:7731 30513</lparam>
<lparam>Address:7732 30514</lparam>
<lparam>Address:7733 30515</lparam>
<lparam>Address:7734 30516</lparam>
<lparam>Address:7735 30517</lparam>
<lparam>Address:7736 30518</lparam>
<lparam>Address:7737 30519</lparam>
<lparam>Address:7738 30520</lparam>
<lparam>Address:7739 30521</lparam>
<lparam>Address:7740 30528</lparam>
<lparam>Address:7741 30529</lparam>
<lparam>Address:7742 30530</lparam>
<lparam>Address:7743 30531</lparam>
<lparam>Address:7744 30532</lparam>
<lparam>Address:7745 30533</lparam>
<lparam>Address:7746 30534</lparam>
<lparam>Address:7747 30535</lparam>
<lparam>Address:7748 30536</lparam>
<lparam>Address:7749 30537</lparam>
<lparam>Address:7750 30544</lparam>
<lparam>Address:7751 30545</lparam>
<lparam>Address:7752 30546</lparam>
<lparam>Address:7753 30547</lparam>
<lparam>Address:7754 30548</lparam>
<lparam>Address:7755 30549</lparam>
<lparam>Address:7756 30550</lparam>
<lparam>Address:7757 30551</lparam>
<lparam>Address:7758 30552</lparam>
<lparam>Address:7759 30553</lparam>
<lparam>Address:7760 30560</lparam>
<lparam>Address:7761 30561</lparam>
<lparam>Address:7762 30562</lparam>
<lparam>Address:7763 30563</lparam>
<lparam>Address:7764 30564</lparam>
<lparam>Address:7765 30565</lparam>
<lparam>Address:7766 30566</lparam>
<lparam>Address:7767 30567</lparam>
<lparam>Address:7768 30568</lparam>
<lparam>Address:7769 30569</lparam>
<lparam>Address:7770 30576</lparam>
<lparam>Address:7771 30577</lparam>
<lparam>Address:7772 30578</lparam>
<lparam>Address:7773 30579</lparam>
<lparam>Address:7774 30580</lparam>
<lparam>Address:7775 30581</lparam>
<lparam>Address:7776 30582</lparam>
<lparam>Address:7777 30583</lparam>
<lparam>Address:7778 30584</lparam>
<lparam>Address:7779 30585</lparam>
<lparam>Address:7780 30592</lparam>
<lparam>Address:7781 30593</lparam>
<lparam>Address:7782 30594</lparam>
<lparam>Address:7783 30595</lparam>
<lparam>Address:7784 30596</lparam>
<lparam>Address:7785 30597</lparam>
<lparam>Address:7786 30598</lparam>
<lparam>Address:7787 30599</lparam>
<lparam>Address:7788 30600</lparam>
<lparam>Address:7789 30601</lparam>
<lparam>Address:7790 30608</lparam>
<lparam>Address:7791 30609</lparam>
<lparam>Address:7792 30610</lparam>
<lparam>Address:7793 30611</lparam>
<lparam>Address:7794 30612</lparam>
<lparam>Address:7795 30613</lparam>
<lparam>Address:7796 30614</lparam>
<lparam>Address:7797 30615</lparam>
<lparam>Address:7798 30616</lparam>
<lparam>Address:7799 30617</lparam>
<lparam>Address:7800 30720</lparam>
<lparam>Address:7801 30721</lparam>
<lparam>Address:7802 30722</lparam>
<lparam>Address:7803 30723</lparam>
<lparam>Address:7804 30724</lparam>
<lparam>Address:7805 30725</lparam>
<lparam>Address:7806 30726</lparam>
<lparam>Address:7807 30727</lparam>
<lparam>Address:7808 30728</lparam>
<lparam>Address:7809 30729</lparam>
<lparam>Address:7810 30736</lparam>
<lparam>Address:7811 30737</lparam>
<lparam>Address:7812 30738</lparam>
<lparam>Address:7813 30739</lparam>
<lparam>Address:7814 30740</lparam>
<lparam>Address:7815 30741</lparam>
<lparam>Address:7816 30742</lparam>
<lparam>Address:7817 30743</lparam>
<lparam>Address:7818 30744</lparam>
<lparam>Address:7819 30745</lparam>
<lparam>Address:7820 30752</lparam>
<lparam>Address:7821 30753</lparam>
<lparam>Address:7822 30754</lparam>
<lparam>Address:7823 30755</lparam>
<lparam>Address:7824 30756</lparam>
<lparam>Address:7825 30757</lparam>
<lparam>Address:7826 30758</lparam>
<lparam>Address:7827 30759</lparam>
<lparam>Address:7828 30760</lparam>
<lparam>Address:7829 30761</lparam>
<lparam>Address:7830 30768</lparam>
<lparam>Address:7831 30769</lparam>
<lparam>Address:7832 30770</lparam>
<lparam>Address:7833 30771</lparam>
<lparam>Address:7834 30772</lparam>
<lparam>Address:7835 30773</lparam>
<lparam>Address:7836 30774</lparam>
<lparam>Address:7837 30775</lparam>
<lparam>Address:7838 30776</lparam>
<lparam>Address:7839 30777</lparam>
<lparam>Address:7840 30784</lparam>
<lparam>Address:7841 30785</lparam>
<lparam>Address:7842 30786</lparam>
<lparam>Address:7843 30787</lparam>
<lparam>Address:7844 30788</lparam>
<lparam>Address:7845 30789</lparam>
<lparam>Address:7846 30790</lparam>
<lparam>Address:7847 30791</lparam>
<lparam>Address:7848 30792</lparam>
<lparam>Address:7849 30793</lparam>
<lparam>Address:7850 30800</lparam>
<lparam>Address:7851 30801</lparam>
<lparam>Address:7852 30802</lparam>
<lparam>Address:7853 30803</lparam>
<lparam>Address:7854 30804</lparam>
<lparam>Address:7855 30805</lparam>
<lparam>Address:7856 30806</lparam>
<lparam>Address:7857 30807</lparam>
<lparam>Address:7858 30808</lparam>
<lparam>Address:7859 30809</lparam>
<lparam>Address:7860 30816</lparam>
<lparam>Address:7861 30817</lparam>
<lparam>Address:7862 30818</lparam>
<lparam>Address:7863 30819</lparam>
<lparam>Address:7864 30820</lparam>
<lparam>Address:7865 30821</lparam>
<lparam>Address:7866 30822</lparam>
<lparam>Address:7867 30823</lparam>
<lparam>Address:7868 30824</lparam>
<lparam>Address:7869 30825</lparam>
<lparam>Address:7870 30832</lparam>
<lparam>Address:7871 30833</lparam>
<lparam>Address:7872 30834</lparam>
<lparam>Address:7873 30835</lparam>
<lparam>Address:7874 30836</lparam>
<lparam>Address:7875 30837</lparam>
<lparam>Address:7876 30838</lparam>
<lparam>Address:7877 30839</lparam>
<lparam>Address:7878 30840</lparam>
<lparam>Address:7879 30841</lparam>
<lparam>Address:7880 30848</lparam>
<lparam>Address:7881 30849</lparam>
<lparam>Address:7882 30850</lparam>
<lparam>Address:7883 30851</lparam>
<lparam>Address:7884 30852</lparam>
<lparam>Address:7885 30853</lparam>
<lparam>Address:7886 30854</lparam>
<lparam>Address:7887 30855</lparam>
<lparam>Address:7888 30856</lparam>
<lparam>Address:7889 30857</lparam>
<lparam>Address:7890 30864</lparam>
<lparam>Address:7891 30865</lparam>
<lparam>Address:7892 30866</lparam>
<lparam>Address:7893 30867</lparam>
<lparam>Address:7894 30868</lparam>
<lparam>Address:7895 30869</lparam>
<lparam>Address:7896 30870</lparam>
<lparam>Address:7897 30871</lparam>
<lparam>Address:7898 30872</lparam>
<lparam>Address:7899 30873</lparam>
<lparam>Address:7900 30976</lparam>
<lparam>Address:7901 30977</lparam>
<lparam>Address:7902 30978</lparam>
<lparam>Address:7903 30979</lparam>
<lparam>Address:7904 30980</lparam>
<lparam>Address:7905 30981</lparam>
<lparam>Address:7906 30982</lparam>
<lparam>Address:7907 30983</lparam>
<lparam>Address:7908 30984</lparam>
<lparam>Address:7909 30985</lparam>
<lparam>Address:7910 30992</lparam>
<lparam>Address:7911 30993</lparam>
<lparam>Address:7912 30994</lparam>
<lparam>Address:7913 30995</lparam>
<lparam>Address:7914 30996</lparam>
<lparam>Address:7915 30997</lparam>
<lparam>Address:7916 30998</lparam>
<lparam>Address:7917 30999</lparam>
<lparam>Address:7918 31000</lparam>
<lparam>Address:7919 31001</lparam>
<lparam>Address:7920 31008</lparam>
<lparam>Address:7921 31009</lparam>
<lparam>Address:7922 31010</lparam>
<lparam>Address:7923 31011</lparam>
<lparam>Address:7924 31012</lparam>
<lparam>Address:7925 31013</lparam>
<lparam>Address:7926 31014</lparam>
<lparam>Address:7927 31015</lparam>
<lparam>Address:7928 31016</lparam>
<lparam>Address:7929 31017</lparam>
<lparam>Address:7930 31024</lparam>
<lparam>Address:7931 31025</lparam>
<lparam>Address:7932 31026</lparam>
<lparam>Address:7933 31027</lparam>
<lparam>Address:7934 31028</lparam>
<lparam>Address:7935 31029</lparam>
<lparam>Address:7936 31030</lparam>
<lparam>Address:7937 31031</lparam>
<lparam>Address:7938 31032</lparam>
<lparam>Address:7939 31033</lparam>
<lparam>Address:7940 31040</lparam>
<lparam>Address:7941 31041</lparam>
<lparam>Address:7942 31042</lparam>
<lparam>Address:7943 31043</lparam>
<lparam>Address:7944 31044</lparam>
<lparam>Address:7945 31045</lparam>
<lparam>Address:7946 31046</lparam>
<lparam>Address:7947 31047</lparam>
<lparam>Address:7948 31048</lparam>
<lparam>Address:7949 31049</lparam>
<lparam>Address:7950 31056</lparam>
<lparam>Address:7951 31057</lparam>
<lparam>Address:7952 31058</lparam>
<lparam>Address:7953 31059</lparam>
<lparam>Address:7954 31060</lparam>
<lparam>Address:7955 31061</lparam>
<lparam>Address:7956 31062</lparam>
<lparam>Address:7957 31063</lparam>
<lparam>Address:7958 31064</lparam>
<lparam>Address:7959 31065</lparam>
<lparam>Address:7960 31072</lparam>
<lparam>Address:7961 31073</lparam>
<lparam>Address:7962 31074</lparam>
<lparam>Address:7963 31075</lparam>
<lparam>Address:7964 31076</lparam>
<lparam>Address:7965 31077</lparam>
<lparam>Address:7966 31078</lparam>
<lparam>Address:7967 31079</lparam>
<lparam>Address:7968 31080</lparam>
<lparam>Address:7969 31081</lparam>
<lparam>Address:7970 31088</lparam>
<lparam>Address:7971 31089</lparam>
<lparam>Address:7972 31090</lparam>
<lparam>Address:7973 31091</lparam>
<lparam>Address:7974 31092</lparam>
<lparam>Address:7975 31093</lparam>
<lparam>Address:7976 31094</lparam>
<lparam>Address:7977 31095</lparam>
<lparam>Address:7978 31096</lparam>
<lparam>Address:7979 31097</lparam>
<lparam>Address:7980 31104</lparam>
<lparam>Address:7981 31105</lparam>
<lparam>Address:7982 31106</lparam>
<lparam>Address:7983 31107</lparam>
<lparam>Address:7984 31108</lparam>
<lparam>Address:7985 31109</lparam>
<lparam>Address:7986 31110</lparam>
<lparam>Address:7987 31111</lparam>
<lparam>Address:7988 31112</lparam>
<lparam>Address:7989 31113</lparam>
<lparam>Address:7990 31120</lparam>
<lparam>Address:7991 31121</lparam>
<lparam>Address:7992 31122</lparam>
<lparam>Address:7993 31123</lparam>
<lparam>Address:7994 31124</lparam>
<lparam>Address:7995 31125</lparam>
<lparam>Address:7996 31126</lparam>
<lparam>Address:7997 31127</lparam>
<lparam>Address:7998 31128</lparam>
<lparam>Address:7999 31129</lparam>
<lparam>Address:8000 28672</lparam>
<lparam>Address:8001 32769</lparam>
<lparam>Address:8002 32770</lparam>
<lparam>Address:8003 32771</lparam>
<lparam>Address:8004 32772</lparam>
<lparam>Address:8005 32773</lparam>
<lparam>Address:8006 32774</lparam>
<lparam>Address:8007 32775</lparam>
<lparam>Address:8008 32776</lparam>
<lparam>Address:8009 32777</lparam>
<lparam>Address:8010 32784</lparam>
<lparam>Address:8011 32785</lparam>
<lparam>Address:8012 32786</lparam>
<lparam>Address:8013 32787</lparam>
<lparam>Address:8014 32788</lparam>
<lparam>Address:8015 32789</lparam>
<lparam>Address:8016 32790</lparam>
<lparam>Address:8017 32791</lparam>
<lparam>Address:8018 32792</lparam>
<lparam>Address:8019 32793</lparam>
<lparam>Address:8020 32800</lparam>
<lparam>Address:8021 32801</lparam>
<lparam>Address:8022 32802</lparam>
<lparam>Address:8023 32803</lparam>
<lparam>Address:8024 32804</lparam>
<lparam>Address:8025 32805</lparam>
<lparam>Address:8026 32806</lparam>
<lparam>Address:8027 32807</lparam>
<lparam>Address:8028 32808</lparam>
<lparam>Address:8029 32809</lparam>
<lparam>Address:8030 32816</lparam>
<lparam>Address:8031 32817</lparam>
<lparam>Address:8032 32818</lparam>
<lparam>Address:8033 32819</lparam>
<lparam>Address:8034 32820</lparam>
<lparam>Address:8035 32821</lparam>
<lparam>Address:8036 32822</lparam>
<lparam>Address:8037 32823</lparam>
<lparam>Address:8038 32824</lparam>
<lparam>Address:8039 32825</lparam>
<lparam>Address:8040 32832</lparam>
<lparam>Address:8041 32833</lparam>
<lparam>Address:8042 32834</lparam>
<lparam>Address:8043 32835</lparam>
<lparam>Address:8044 32836</lparam>
<lparam>Address:8045 32837</lparam>
<lparam>Address:8046 32838</lparam>
<lparam>Address:8047 32839</lparam>
<lparam>Address:8048 32840</lparam>
<lparam>Address:8049 32841</lparam>
<lparam>Address:8050 32848</lparam>
<lparam>Address:8051 32849</lparam>
<lparam>Address:8052 32850</lparam>
<lparam>Address:8053 32851</lparam>
<lparam>Address:8054 32852</lparam>
<lparam>Address:8055 32853</lparam>
<lparam>Address:8056 32854</lparam>
<lparam>Address:8057 32855</lparam>
<lparam>Address:8058 32856</lparam>
<lparam>Address:8059 32857</lparam>
<lparam>Address:8060 32864</lparam>
<lparam>Address:8061 32865</lparam>
<lparam>Address:8062 32866</lparam>
<lparam>Address:8063 32867</lparam>
<lparam>Address:8064 32868</lparam>
<lparam>Address:8065 32869</lparam>
<lparam>Address:8066 32870</lparam>
<lparam>Address:8067 32871</lparam>
<lparam>Address:8068 32872</lparam>
<lparam>Address:8069 32873</lparam>
<lparam>Address:8070 32880</lparam>
<lparam>Address:8071 32881</lparam>
<lparam>Address:8072 32882</lparam>
<lparam>Address:8073 32883</lparam>
<lparam>Address:8074 32884</lparam>
<lparam>Address:8075 32885</lparam>
<lparam>Address:8076 32886</lparam>
<lparam>Address:8077 32887</lparam>
<lparam>Address:8078 32888</lparam>
<lparam>Address:8079 32889</lparam>
<lparam>Address:8080 32896</lparam>
<lparam>Address:8081 32897</lparam>
<lparam>Address:8082 32898</lparam>
<lparam>Address:8083 32899</lparam>
<lparam>Address:8084 32900</lparam>
<lparam>Address:8085 32901</lparam>
<lparam>Address:8086 32902</lparam>
<lparam>Address:8087 32903</lparam>
<lparam>Address:8088 32904</lparam>
<lparam>Address:8089 32905</lparam>
<lparam>Address:8090 32912</lparam>
<lparam>Address:8091 32913</lparam>
<lparam>Address:8092 32914</lparam>
<lparam>Address:8093 32915</lparam>
<lparam>Address:8094 32916</lparam>
<lparam>Address:8095 32917</lparam>
<lparam>Address:8096 32918</lparam>
<lparam>Address:8097 32919</lparam>
<lparam>Address:8098 32920</lparam>
<lparam>Address:8099 32921</lparam>
<lparam>Address:8100 33024</lparam>
<lparam>Address:8101 33025</lparam>
<lparam>Address:8102 33026</lparam>
<lparam>Address:8103 33027</lparam>
<lparam>Address:8104 33028</lparam>
<lparam>Address:8105 33029</lparam>
<lparam>Address:8106 33030</lparam>
<lparam>Address:8107 33031</lparam>
<lparam>Address:8108 33032</lparam>
<lparam>Address:8109 33033</lparam>
<lparam>Address:8110 33040</lparam>
<lparam>Address:8111 33041</lparam>
<lparam>Address:8112 33042</lparam>
<lparam>Address:8113 33043</lparam>
<lparam>Address:8114 33044</lparam>
<lparam>Address:8115 33045</lparam>
<lparam>Address:8116 33046</lparam>
<lparam>Address:8117 33047</lparam>
<lparam>Address:8118 33048</lparam>
<lparam>Address:8119 33049</lparam>
<lparam>Address:8120 33056</lparam>
<lparam>Address:8121 33057</lparam>
<lparam>Address:8122 33058</lparam>
<lparam>Address:8123 33059</lparam>
<lparam>Address:8124 33060</lparam>
<lparam>Address:8125 33061</lparam>
<lparam>Address:8126 33062</lparam>
<lparam>Address:8127 33063</lparam>
<lparam>Address:8128 33064</lparam>
<lparam>Address:8129 33065</lparam>
<lparam>Address:8130 33072</lparam>
<lparam>Address:8131 33073</lparam>
<lparam>Address:8132 33074</lparam>
<lparam>Address:8133 33075</lparam>
<lparam>Address:8134 33076</lparam>
<lparam>Address:8135 33077</lparam>
<lparam>Address:8136 33078</lparam>
<lparam>Address:8137 33079</lparam>
<lparam>Address:8138 33080</lparam>
<lparam>Address:8139 33081</lparam>
<lparam>Address:8140 33088</lparam>
<lparam>Address:8141 33089</lparam>
<lparam>Address:8142 33090</lparam>
<lparam>Address:8143 33091</lparam>
<lparam>Address:8144 33092</lparam>
<lparam>Address:8145 33093</lparam>
<lparam>Address:8146 33094</lparam>
<lparam>Address:8147 33095</lparam>
<lparam>Address:8148 33096</lparam>
<lparam>Address:8149 33097</lparam>
<lparam>Address:8150 33104</lparam>
<lparam>Address:8151 33105</lparam>
<lparam>Address:8152 33106</lparam>
<lparam>Address:8153 33107</lparam>
<lparam>Address:8154 33108</lparam>
<lparam>Address:8155 33109</lparam>
<lparam>Address:8156 33110</lparam>
<lparam>Address:8157 33111</lparam>
<lparam>Address:8158 33112</lparam>
<lparam>Address:8159 33113</lparam>
<lparam>Address:8160 33120</lparam>
<lparam>Address:8161 33121</lparam>
<lparam>Address:8162 33122</lparam>
<lparam>Address:8163 33123</lparam>
<lparam>Address:8164 33124</lparam>
<lparam>Address:8165 33125</lparam>
<lparam>Address:8166 33126</lparam>
<lparam>Address:8167 33127</lparam>
<lparam>Address:8168 33128</lparam>
<lparam>Address:8169 33129</lparam>
<lparam>Address:8170 33136</lparam>
<lparam>Address:8171 33137</lparam>
<lparam>Address:8172 33138</lparam>
<lparam>Address:8173 33139</lparam>
<lparam>Address:8174 33140</lparam>
<lparam>Address:8175 33141</lparam>
<lparam>Address:8176 33142</lparam>
<lparam>Address:8177 33143</lparam>
<lparam>Address:8178 33144</lparam>
<lparam>Address:8179 33145</lparam>
<lparam>Address:8180 33152</lparam>
<lparam>Address:8181 33153</lparam>
<lparam>Address:8182 33154</lparam>
<lparam>Address:8183 33155</lparam>
<lparam>Address:8184 33156</lparam>
<lparam>Address:8185 33157</lparam>
<lparam>Address:8186 33158</lparam>
<lparam>Address:8187 33159</lparam>
<lparam>Address:8188 33160</lparam>
<lparam>Address:8189 33161</lparam>
<lparam>Address:8190 33168</lparam>
<lparam>Address:8191 33169</lparam>
<lparam>Address:8192 33170</lparam>
<lparam>Address:8193 33171</lparam>
<lparam>Address:8194 33172</lparam>
<lparam>Address:8195 33173</lparam>
<lparam>Address:8196 33174</lparam>
<lparam>Address:8197 33175</lparam>
<lparam>Address:8198 33176</lparam>
<lparam>Address:8199 33177</lparam>
<lparam>Address:8200 33280</lparam>
<lparam>Address:8201 33281</lparam>
<lparam>Address:8202 33282</lparam>
<lparam>Address:8203 33283</lparam>
<lparam>Address:8204 33284</lparam>
<lparam>Address:8205 33285</lparam>
<lparam>Address:8206 33286</lparam>
<lparam>Address:8207 33287</lparam>
<lparam>Address:8208 33288</lparam>
<lparam>Address:8209 33289</lparam>
<lparam>Address:8210 33296</lparam>
<lparam>Address:8211 33297</lparam>
<lparam>Address:8212 33298</lparam>
<lparam>Address:8213 33299</lparam>
<lparam>Address:8214 33300</lparam>
<lparam>Address:8215 33301</lparam>
<lparam>Address:8216 33302</lparam>
<lparam>Address:8217 33303</lparam>
<lparam>Address:8218 33304</lparam>
<lparam>Address:8219 33305</lparam>
<lparam>Address:8220 33312</lparam>
<lparam>Address:8221 33313</lparam>
<lparam>Address:8222 33314</lparam>
<lparam>Address:8223 33315</lparam>
<lparam>Address:8224 33316</lparam>
<lparam>Address:8225 33317</lparam>
<lparam>Address:8226 33318</lparam>
<lparam>Address:8227 33319</lparam>
<lparam>Address:8228 33320</lparam>
<lparam>Address:8229 33321</lparam>
<lparam>Address:8230 33328</lparam>
<lparam>Address:8231 33329</lparam>
<lparam>Address:8232 33330</lparam>
<lparam>Address:8233 33331</lparam>
<lparam>Address:8234 33332</lparam>
<lparam>Address:8235 33333</lparam>
<lparam>Address:8236 33334</lparam>
<lparam>Address:8237 33335</lparam>
<lparam>Address:8238 33336</lparam>
<lparam>Address:8239 33337</lparam>
<lparam>Address:8240 33344</lparam>
<lparam>Address:8241 33345</lparam>
<lparam>Address:8242 33346</lparam>
<lparam>Address:8243 33347</lparam>
<lparam>Address:8244 33348</lparam>
<lparam>Address:8245 33349</lparam>
<lparam>Address:8246 33350</lparam>
<lparam>Address:8247 33351</lparam>
<lparam>Address:8248 33352</lparam>
<lparam>Address:8249 33353</lparam>
<lparam>Address:8250 33360</lparam>
<lparam>Address:8251 33361</lparam>
<lparam>Address:8252 33362</lparam>
<lparam>Address:8253 33363</lparam>
<lparam>Address:8254 33364</lparam>
<lparam>Address:8255 33365</lparam>
<lparam>Address:8256 33366</lparam>
<lparam>Address:8257 33367</lparam>
<lparam>Address:8258 33368</lparam>
<lparam>Address:8259 33369</lparam>
<lparam>Address:8260 33376</lparam>
<lparam>Address:8261 33377</lparam>
<lparam>Address:8262 33378</lparam>
<lparam>Address:8263 33379</lparam>
<lparam>Address:8264 33380</lparam>
<lparam>Address:8265 33381</lparam>
<lparam>Address:8266 33382</lparam>
<lparam>Address:8267 33383</lparam>
<lparam>Address:8268 33384</lparam>
<lparam>Address:8269 33385</lparam>
<lparam>Address:8270 33392</lparam>
<lparam>Address:8271 33393</lparam>
<lparam>Address:8272 33394</lparam>
<lparam>Address:8273 33395</lparam>
<lparam>Address:8274 33396</lparam>
<lparam>Address:8275 33397</lparam>
<lparam>Address:8276 33398</lparam>
<lparam>Address:8277 33399</lparam>
<lparam>Address:8278 33400</lparam>
<lparam>Address:8279 33401</lparam>
<lparam>Address:8280 33408</lparam>
<lparam>Address:8281 33409</lparam>
<lparam>Address:8282 33410</lparam>
<lparam>Address:8283 33411</lparam>
<lparam>Address:8284 33412</lparam>
<lparam>Address:8285 33413</lparam>
<lparam>Address:8286 33414</lparam>
<lparam>Address:8287 33415</lparam>
<lparam>Address:8288 33416</lparam>
<lparam>Address:8289 33417</lparam>
<lparam>Address:8290 33424</lparam>
<lparam>Address:8291 33425</lparam>
<lparam>Address:8292 33426</lparam>
<lparam>Address:8293 33427</lparam>
<lparam>Address:8294 33428</lparam>
<lparam>Address:8295 33429</lparam>
<lparam>Address:8296 33430</lparam>
<lparam>Address:8297 33431</lparam>
<lparam>Address:8298 33432</lparam>
<lparam>Address:8299 33433</lparam>
<lparam>Address:8300 33536</lparam>
<lparam>Address:8301 33537</lparam>
<lparam>Address:8302 33538</lparam>
<lparam>Address:8303 33539</lparam>
<lparam>Address:8304 33540</lparam>
<lparam>Address:8305 33541</lparam>
<lparam>Address:8306 33542</lparam>
<lparam>Address:8307 33543</lparam>
<lparam>Address:8308 33544</lparam>
<lparam>Address:8309 33545</lparam>
<lparam>Address:8310 33552</lparam>
<lparam>Address:8311 33553</lparam>
<lparam>Address:8312 33554</lparam>
<lparam>Address:8313 33555</lparam>
<lparam>Address:8314 33556</lparam>
<lparam>Address:8315 33557</lparam>
<lparam>Address:8316 33558</lparam>
<lparam>Address:8317 33559</lparam>
<lparam>Address:8318 33560</lparam>
<lparam>Address:8319 33561</lparam>
<lparam>Address:8320 33568</lparam>
<lparam>Address:8321 33569</lparam>
<lparam>Address:8322 33570</lparam>
<lparam>Address:8323 33571</lparam>
<lparam>Address:8324 33572</lparam>
<lparam>Address:8325 33573</lparam>
<lparam>Address:8326 33574</lparam>
<lparam>Address:8327 33575</lparam>
<lparam>Address:8328 33576</lparam>
<lparam>Address:8329 33577</lparam>
<lparam>Address:8330 33584</lparam>
<lparam>Address:8331 33585</lparam>
<lparam>Address:8332 33586</lparam>
<lparam>Address:8333 33587</lparam>
<lparam>Address:8334 33588</lparam>
<lparam>Address:8335 33589</lparam>
<lparam>Address:8336 33590</lparam>
<lparam>Address:8337 33591</lparam>
<lparam>Address:8338 33592</lparam>
<lparam>Address:8339 33593</lparam>
<lparam>Address:8340 33600</lparam>
<lparam>Address:8341 33601</lparam>
<lparam>Address:8342 33602</lparam>
<lparam>Address:8343 33603</lparam>
<lparam>Address:8344 33604</lparam>
<lparam>Address:8345 33605</lparam>
<lparam>Address:8346 33606</lparam>
<lparam>Address:8347 33607</lparam>
<lparam>Address:8348 33608</lparam>
<lparam>Address:8349 33609</lparam>
<lparam>Address:8350 33616</lparam>
<lparam>Address:8351 33617</lparam>
<lparam>Address:8352 33618</lparam>
<lparam>Address:8353 33619</lparam>
<lparam>Address:8354 33620</lparam>
<lparam>Address:8355 33621</lparam>
<lparam>Address:8356 33622</lparam>
<lparam>Address:8357 33623</lparam>
<lparam>Address:8358 33624</lparam>
<lparam>Address:8359 33625</lparam>
<lparam>Address:8360 33632</lparam>
<lparam>Address:8361 33633</lparam>
<lparam>Address:8362 33634</lparam>
<lparam>Address:8363 33635</lparam>
<lparam>Address:8364 33636</lparam>
<lparam>Address:8365 33637</lparam>
<lparam>Address:8366 33638</lparam>
<lparam>Address:8367 33639</lparam>
<lparam>Address:8368 33640</lparam>
<lparam>Address:8369 33641</lparam>
<lparam>Address:8370 33648</lparam>
<lparam>Address:8371 33649</lparam>
<lparam>Address:8372 33650</lparam>
<lparam>Address:8373 33651</lparam>
<lparam>Address:8374 33652</lparam>
<lparam>Address:8375 33653</lparam>
<lparam>Address:8376 33654</lparam>
<lparam>Address:8377 33655</lparam>
<lparam>Address:8378 33656</lparam>
<lparam>Address:8379 33657</lparam>
<lparam>Address:8380 33664</lparam>
<lparam>Address:8381 33665</lparam>
<lparam>Address:8382 33666</lparam>
<lparam>Address:8383 33667</lparam>
<lparam>Address:8384 33668</lparam>
<lparam>Address:8385 33669</lparam>
<lparam>Address:8386 33670</lparam>
<lparam>Address:8387 33671</lparam>
<lparam>Address:8388 33672</lparam>
<lparam>Address:8389 33673</lparam>
<lparam>Address:8390 33680</lparam>
<lparam>Address:8391 33681</lparam>
<lparam>Address:8392 33682</lparam>
<lparam>Address:8393 33683</lparam>
<lparam>Address:8394 33684</lparam>
<lparam>Address:8395 33685</lparam>
<lparam>Address:8396 33686</lparam>
<lparam>Address:8397 33687</lparam>
<lparam>Address:8398 33688</lparam>
<lparam>Address:8399 33689</lparam>
<lparam>Address:8400 33792</lparam>
<lparam>Address:8401 33793</lparam>
<lparam>Address:8402 33794</lparam>
<lparam>Address:8403 33795</lparam>
<lparam>Address:8404 33796</lparam>
<lparam>Address:8405 33797</lparam>
<lparam>Address:8406 33798</lparam>
<lparam>Address:8407 33799</lparam>
<lparam>Address:8408 33800</lparam>
<lparam>Address:8409 33801</lparam>
<lparam>Address:8410 33808</lparam>
<lparam>Address:8411 33809</lparam>
<lparam>Address:8412 33810</lparam>
<lparam>Address:8413 33811</lparam>
<lparam>Address:8414 33812</lparam>
<lparam>Address:8415 33813</lparam>
<lparam>Address:8416 33814</lparam>
<lparam>Address:8417 33815</lparam>
<lparam>Address:8418 33816</lparam>
<lparam>Address:8419 33817</lparam>
<lparam>Address:8420 33824</lparam>
<lparam>Address:8421 33825</lparam>
<lparam>Address:8422 33826</lparam>
<lparam>Address:8423 33827</lparam>
<lparam>Address:8424 33828</lparam>
<lparam>Address:8425 33829</lparam>
<lparam>Address:8426 33830</lparam>
<lparam>Address:8427 33831</lparam>
<lparam>Address:8428 33832</lparam>
<lparam>Address:8429 33833</lparam>
<lparam>Address:8430 33840</lparam>
<lparam>Address:8431 33841</lparam>
<lparam>Address:8432 33842</lparam>
<lparam>Address:8433 33843</lparam>
<lparam>Address:8434 33844</lparam>
<lparam>Address:8435 33845</lparam>
<lparam>Address:8436 33846</lparam>
<lparam>Address:8437 33847</lparam>
<lparam>Address:8438 33848</lparam>
<lparam>Address:8439 33849</lparam>
<lparam>Address:8440 33856</lparam>
<lparam>Address:8441 33857</lparam>
<lparam>Address:8442 33858</lparam>
<lparam>Address:8443 33859</lparam>
<lparam>Address:8444 33860</lparam>
<lparam>Address:8445 33861</lparam>
<lparam>Address:8446 33862</lparam>
<lparam>Address:8447 33863</lparam>
<lparam>Address:8448 33864</lparam>
<lparam>Address:8449 33865</lparam>
<lparam>Address:8450 33872</lparam>
<lparam>Address:8451 33873</lparam>
<lparam>Address:8452 33874</lparam>
<lparam>Address:8453 33875</lparam>
<lparam>Address:8454 33876</lparam>
<lparam>Address:8455 33877</lparam>
<lparam>Address:8456 33878</lparam>
<lparam>Address:8457 33879</lparam>
<lparam>Address:8458 33880</lparam>
<lparam>Address:8459 33881</lparam>
<lparam>Address:8460 33888</lparam>
<lparam>Address:8461 33889</lparam>
<lparam>Address:8462 33890</lparam>
<lparam>Address:8463 33891</lparam>
<lparam>Address:8464 33892</lparam>
<lparam>Address:8465 33893</lparam>
<lparam>Address:8466 33894</lparam>
<lparam>Address:8467 33895</lparam>
<lparam>Address:8468 33896</lparam>
<lparam>Address:8469 33897</lparam>
<lparam>Address:8470 33904</lparam>
<lparam>Address:8471 33905</lparam>
<lparam>Address:8472 33906</lparam>
<lparam>Address:8473 33907</lparam>
<lparam>Address:8474 33908</lparam>
<lparam>Address:8475 33909</lparam>
<lparam>Address:8476 33910</lparam>
<lparam>Address:8477 33911</lparam>
<lparam>Address:8478 33912</lparam>
<lparam>Address:8479 33913</lparam>
<lparam>Address:8480 33920</lparam>
<lparam>Address:8481 33921</lparam>
<lparam>Address:8482 33922</lparam>
<lparam>Address:8483 33923</lparam>
<lparam>Address:8484 33924</lparam>
<lparam>Address:8485 33925</lparam>
<lparam>Address:8486 33926</lparam>
<lparam>Address:8487 33927</lparam>
<lparam>Address:8488 33928</lparam>
<lparam>Address:8489 33929</lparam>
<lparam>Address:8490 33936</lparam>
<lparam>Address:8491 33937</lparam>
<lparam>Address:8492 33938</lparam>
<lparam>Address:8493 33939</lparam>
<lparam>Address:8494 33940</lparam>
<lparam>Address:8495 33941</lparam>
<lparam>Address:8496 33942</lparam>
<lparam>Address:8497 33943</lparam>
<lparam>Address:8498 33944</lparam>
<lparam>Address:8499 33945</lparam>
<lparam>Address:8500 34048</lparam>
<lparam>Address:8501 34049</lparam>
<lparam>Address:8502 34050</lparam>
<lparam>Address:8503 34051</lparam>
<lparam>Address:8504 34052</lparam>
<lparam>Address:8505 34053</lparam>
<lparam>Address:8506 34054</lparam>
<lparam>Address:8507 34055</lparam>
<lparam>Address:8508 34056</lparam>
<lparam>Address:8509 34057</lparam>
<lparam>Address:8510 34064</lparam>
<lparam>Address:8511 34065</lparam>
<lparam>Address:8512 34066</lparam>
<lparam>Address:8513 34067</lparam>
<lparam>Address:8514 34068</lparam>
<lparam>Address:8515 34069</lparam>
<lparam>Address:8516 34070</lparam>
<lparam>Address:8517 34071</lparam>
<lparam>Address:8518 34072</lparam>
<lparam>Address:8519 34073</lparam>
<lparam>Address:8520 34080</lparam>
<lparam>Address:8521 34081</lparam>
<lparam>Address:8522 34082</lparam>
<lparam>Address:8523 34083</lparam>
<lparam>Address:8524 34084</lparam>
<lparam>Address:8525 34085</lparam>
<lparam>Address:8526 34086</lparam>
<lparam>Address:8527 34087</lparam>
<lparam>Address:8528 34088</lparam>
<lparam>Address:8529 34089</lparam>
<lparam>Address:8530 34096</lparam>
<lparam>Address:8531 34097</lparam>
<lparam>Address:8532 34098</lparam>
<lparam>Address:8533 34099</lparam>
<lparam>Address:8534 34100</lparam>
<lparam>Address:8535 34101</lparam>
<lparam>Address:8536 34102</lparam>
<lparam>Address:8537 34103</lparam>
<lparam>Address:8538 34104</lparam>
<lparam>Address:8539 34105</lparam>
<lparam>Address:8540 34112</lparam>
<lparam>Address:8541 34113</lparam>
<lparam>Address:8542 34114</lparam>
<lparam>Address:8543 34115</lparam>
<lparam>Address:8544 34116</lparam>
<lparam>Address:8545 34117</lparam>
<lparam>Address:8546 34118</lparam>
<lparam>Address:8547 34119</lparam>
<lparam>Address:8548 34120</lparam>
<lparam>Address:8549 34121</lparam>
<lparam>Address:8550 34128</lparam>
<lparam>Address:8551 34129</lparam>
<lparam>Address:8552 34130</lparam>
<lparam>Address:8553 34131</lparam>
<lparam>Address:8554 34132</lparam>
<lparam>Address:8555 34133</lparam>
<lparam>Address:8556 34134</lparam>
<lparam>Address:8557 34135</lparam>
<lparam>Address:8558 34136</lparam>
<lparam>Address:8559 34137</lparam>
<lparam>Address:8560 34144</lparam>
<lparam>Address:8561 34145</lparam>
<lparam>Address:8562 34146</lparam>
<lparam>Address:8563 34147</lparam>
<lparam>Address:8564 34148</lparam>
<lparam>Address:8565 34149</lparam>
<lparam>Address:8566 34150</lparam>
<lparam>Address:8567 34151</lparam>
<lparam>Address:8568 34152</lparam>
<lparam>Address:8569 34153</lparam>
<lparam>Address:8570 34160</lparam>
<lparam>Address:8571 34161</lparam>
<lparam>Address:8572 34162</lparam>
<lparam>Address:8573 34163</lparam>
<lparam>Address:8574 34164</lparam>
<lparam>Address:8575 34165</lparam>
<lparam>Address:8576 34166</lparam>
<lparam>Address:8577 34167</lparam>
<lparam>Address:8578 34168</lparam>
<lparam>Address:8579 34169</lparam>
<lparam>Address:8580 34176</lparam>
<lparam>Address:8581 34177</lparam>
<lparam>Address:8582 34178</lparam>
<lparam>Address:8583 34179</lparam>
<lparam>Address:8584 34180</lparam>
<lparam>Address:8585 34181</lparam>
<lparam>Address:8586 34182</lparam>
<lparam>Address:8587 34183</lparam>
<lparam>Address:8588 34184</lparam>
<lparam>Address:8589 34185</lparam>
<lparam>Address:8590 34192</lparam>
<lparam>Address:8591 34193</lparam>
<lparam>Address:8592 34194</lparam>
<lparam>Address:8593 34195</lparam>
<lparam>Address:8594 34196</lparam>
<lparam>Address:8595 34197</lparam>
<lparam>Address:8596 34198</lparam>
<lparam>Address:8597 34199</lparam>
<lparam>Address:8598 34200</lparam>
<lparam>Address:8599 34201</lparam>
<lparam>Address:8600 34304</lparam>
<lparam>Address:8601 34305</lparam>
<lparam>Address:8602 34306</lparam>
<lparam>Address:8603 34307</lparam>
<lparam>Address:8604 34308</lparam>
<lparam>Address:8605 34309</lparam>
<lparam>Address:8606 34310</lparam>
<lparam>Address:8607 34311</lparam>
<lparam>Address:8608 34312</lparam>
<lparam>Address:8609 34313</lparam>
<lparam>Address:8610 34320</lparam>
<lparam>Address:8611 34321</lparam>
<lparam>Address:8612 34322</lparam>
<lparam>Address:8613 34323</lparam>
<lparam>Address:8614 34324</lparam>
<lparam>Address:8615 34325</lparam>
<lparam>Address:8616 34326</lparam>
<lparam>Address:8617 34327</lparam>
<lparam>Address:8618 34328</lparam>
<lparam>Address:8619 34329</lparam>
<lparam>Address:8620 34336</lparam>
<lparam>Address:8621 34337</lparam>
<lparam>Address:8622 34338</lparam>
<lparam>Address:8623 34339</lparam>
<lparam>Address:8624 34340</lparam>
<lparam>Address:8625 34341</lparam>
<lparam>Address:8626 34342</lparam>
<lparam>Address:8627 34343</lparam>
<lparam>Address:8628 34344</lparam>
<lparam>Address:8629 34345</lparam>
<lparam>Address:8630 34352</lparam>
<lparam>Address:8631 34353</lparam>
<lparam>Address:8632 34354</lparam>
<lparam>Address:8633 34355</lparam>
<lparam>Address:8634 34356</lparam>
<lparam>Address:8635 34357</lparam>
<lparam>Address:8636 34358</lparam>
<lparam>Address:8637 34359</lparam>
<lparam>Address:8638 34360</lparam>
<lparam>Address:8639 34361</lparam>
<lparam>Address:8640 34368</lparam>
<lparam>Address:8641 34369</lparam>
<lparam>Address:8642 34370</lparam>
<lparam>Address:8643 34371</lparam>
<lparam>Address:8644 34372</lparam>
<lparam>Address:8645 34373</lparam>
<lparam>Address:8646 34374</lparam>
<lparam>Address:8647 34375</lparam>
<lparam>Address:8648 34376</lparam>
<lparam>Address:8649 34377</lparam>
<lparam>Address:8650 34384</lparam>
<lparam>Address:8651 34385</lparam>
<lparam>Address:8652 34386</lparam>
<lparam>Address:8653 34387</lparam>
<lparam>Address:8654 34388</lparam>
<lparam>Address:8655 34389</lparam>
<lparam>Address:8656 34390</lparam>
<lparam>Address:8657 34391</lparam>
<lparam>Address:8658 34392</lparam>
<lparam>Address:8659 34393</lparam>
<lparam>Address:8660 34400</lparam>
<lparam>Address:8661 34401</lparam>
<lparam>Address:8662 34402</lparam>
<lparam>Address:8663 34403</lparam>
<lparam>Address:8664 34404</lparam>
<lparam>Address:8665 34405</lparam>
<lparam>Address:8666 34406</lparam>
<lparam>Address:8667 34407</lparam>
<lparam>Address:8668 34408</lparam>
<lparam>Address:8669 34409</lparam>
<lparam>Address:8670 34416</lparam>
<lparam>Address:8671 34417</lparam>
<lparam>Address:8672 34418</lparam>
<lparam>Address:8673 34419</lparam>
<lparam>Address:8674 34420</lparam>
<lparam>Address:8675 34421</lparam>
<lparam>Address:8676 34422</lparam>
<lparam>Address:8677 34423</lparam>
<lparam>Address:8678 34424</lparam>
<lparam>Address:8679 34425</lparam>
<lparam>Address:8680 34432</lparam>
<lparam>Address:8681 34433</lparam>
<lparam>Address:8682 34434</lparam>
<lparam>Address:8683 34435</lparam>
<lparam>Address:8684 34436</lparam>
<lparam>Address:8685 34437</lparam>
<lparam>Address:8686 34438</lparam>
<lparam>Address:8687 34439</lparam>
<lparam>Address:8688 34440</lparam>
<lparam>Address:8689 34441</lparam>
<lparam>Address:8690 34448</lparam>
<lparam>Address:8691 34449</lparam>
<lparam>Address:8692 34450</lparam>
<lparam>Address:8693 34451</lparam>
<lparam>Address:8694 34452</lparam>
<lparam>Address:8695 34453</lparam>
<lparam>Address:8696 34454</lparam>
<lparam>Address:8697 34455</lparam>
<lparam>Address:8698 34456</lparam>
<lparam>Address:8699 34457</lparam>
<lparam>Address:8700 34560</lparam>
<lparam>Address:8701 34561</lparam>
<lparam>Address:8702 34562</lparam>
<lparam>Address:8703 34563</lparam>
<lparam>Address:8704 34564</lparam>
<lparam>Address:8705 34565</lparam>
<lparam>Address:8706 34566</lparam>
<lparam>Address:8707 34567</lparam>
<lparam>Address:8708 34568</lparam>
<lparam>Address:8709 34569</lparam>
<lparam>Address:8710 34576</lparam>
<lparam>Address:8711 34577</lparam>
<lparam>Address:8712 34578</lparam>
<lparam>Address:8713 34579</lparam>
<lparam>Address:8714 34580</lparam>
<lparam>Address:8715 34581</lparam>
<lparam>Address:8716 34582</lparam>
<lparam>Address:8717 34583</lparam>
<lparam>Address:8718 34584</lparam>
<lparam>Address:8719 34585</lparam>
<lparam>Address:8720 34592</lparam>
<lparam>Address:8721 34593</lparam>
<lparam>Address:8722 34594</lparam>
<lparam>Address:8723 34595</lparam>
<lparam>Address:8724 34596</lparam>
<lparam>Address:8725 34597</lparam>
<lparam>Address:8726 34598</lparam>
<lparam>Address:8727 34599</lparam>
<lparam>Address:8728 34600</lparam>
<lparam>Address:8729 34601</lparam>
<lparam>Address:8730 34608</lparam>
<lparam>Address:8731 34609</lparam>
<lparam>Address:8732 34610</lparam>
<lparam>Address:8733 34611</lparam>
<lparam>Address:8734 34612</lparam>
<lparam>Address:8735 34613</lparam>
<lparam>Address:8736 34614</lparam>
<lparam>Address:8737 34615</lparam>
<lparam>Address:8738 34616</lparam>
<lparam>Address:8739 34617</lparam>
<lparam>Address:8740 34624</lparam>
<lparam>Address:8741 34625</lparam>
<lparam>Address:8742 34626</lparam>
<lparam>Address:8743 34627</lparam>
<lparam>Address:8744 34628</lparam>
<lparam>Address:8745 34629</lparam>
<lparam>Address:8746 34630</lparam>
<lparam>Address:8747 34631</lparam>
<lparam>Address:8748 34632</lparam>
<lparam>Address:8749 34633</lparam>
<lparam>Address:8750 34640</lparam>
<lparam>Address:8751 34641</lparam>
<lparam>Address:8752 34642</lparam>
<lparam>Address:8753 34643</lparam>
<lparam>Address:8754 34644</lparam>
<lparam>Address:8755 34645</lparam>
<lparam>Address:8756 34646</lparam>
<lparam>Address:8757 34647</lparam>
<lparam>Address:8758 34648</lparam>
<lparam>Address:8759 34649</lparam>
<lparam>Address:8760 34656</lparam>
<lparam>Address:8761 34657</lparam>
<lparam>Address:8762 34658</lparam>
<lparam>Address:8763 34659</lparam>
<lparam>Address:8764 34660</lparam>
<lparam>Address:8765 34661</lparam>
<lparam>Address:8766 34662</lparam>
<lparam>Address:8767 34663</lparam>
<lparam>Address:8768 34664</lparam>
<lparam>Address:8769 34665</lparam>
<lparam>Address:8770 34672</lparam>
<lparam>Address:8771 34673</lparam>
<lparam>Address:8772 34674</lparam>
<lparam>Address:8773 34675</lparam>
<lparam>Address:8774 34676</lparam>
<lparam>Address:8775 34677</lparam>
<lparam>Address:8776 34678</lparam>
<lparam>Address:8777 34679</lparam>
<lparam>Address:8778 34680</lparam>
<lparam>Address:8779 34681</lparam>
<lparam>Address:8780 34688</lparam>
<lparam>Address:8781 34689</lparam>
<lparam>Address:8782 34690</lparam>
<lparam>Address:8783 34691</lparam>
<lparam>Address:8784 34692</lparam>
<lparam>Address:8785 34693</lparam>
<lparam>Address:8786 34694</lparam>
<lparam>Address:8787 34695</lparam>
<lparam>Address:8788 34696</lparam>
<lparam>Address:8789 34697</lparam>
<lparam>Address:8790 34704</lparam>
<lparam>Address:8791 34705</lparam>
<lparam>Address:8792 34706</lparam>
<lparam>Address:8793 34707</lparam>
<lparam>Address:8794 34708</lparam>
<lparam>Address:8795 34709</lparam>
<lparam>Address:8796 34710</lparam>
<lparam>Address:8797 34711</lparam>
<lparam>Address:8798 34712</lparam>
<lparam>Address:8799 34713</lparam>
<lparam>Address:8800 34816</lparam>
<lparam>Address:8801 34817</lparam>
<lparam>Address:8802 34818</lparam>
<lparam>Address:8803 34819</lparam>
<lparam>Address:8804 34820</lparam>
<lparam>Address:8805 34821</lparam>
<lparam>Address:8806 34822</lparam>
<lparam>Address:8807 34823</lparam>
<lparam>Address:8808 34824</lparam>
<lparam>Address:8809 34825</lparam>
<lparam>Address:8810 34832</lparam>
<lparam>Address:8811 34833</lparam>
<lparam>Address:8812 34834</lparam>
<lparam>Address:8813 34835</lparam>
<lparam>Address:8814 34836</lparam>
<lparam>Address:8815 34837</lparam>
<lparam>Address:8816 34838</lparam>
<lparam>Address:8817 34839</lparam>
<lparam>Address:8818 34840</lparam>
<lparam>Address:8819 34841</lparam>
<lparam>Address:8820 34848</lparam>
<lparam>Address:8821 34849</lparam>
<lparam>Address:8822 34850</lparam>
<lparam>Address:8823 34851</lparam>
<lparam>Address:8824 34852</lparam>
<lparam>Address:8825 34853</lparam>
<lparam>Address:8826 34854</lparam>
<lparam>Address:8827 34855</lparam>
<lparam>Address:8828 34856</lparam>
<lparam>Address:8829 34857</lparam>
<lparam>Address:8830 34864</lparam>
<lparam>Address:8831 34865</lparam>
<lparam>Address:8832 34866</lparam>
<lparam>Address:8833 34867</lparam>
<lparam>Address:8834 34868</lparam>
<lparam>Address:8835 34869</lparam>
<lparam>Address:8836 34870</lparam>
<lparam>Address:8837 34871</lparam>
<lparam>Address:8838 34872</lparam>
<lparam>Address:8839 34873</lparam>
<lparam>Address:8840 34880</lparam>
<lparam>Address:8841 34881</lparam>
<lparam>Address:8842 34882</lparam>
<lparam>Address:8843 34883</lparam>
<lparam>Address:8844 34884</lparam>
<lparam>Address:8845 34885</lparam>
<lparam>Address:8846 34886</lparam>
<lparam>Address:8847 34887</lparam>
<lparam>Address:8848 34888</lparam>
<lparam>Address:8849 34889</lparam>
<lparam>Address:8850 34896</lparam>
<lparam>Address:8851 34897</lparam>
<lparam>Address:8852 34898</lparam>
<lparam>Address:8853 34899</lparam>
<lparam>Address:8854 34900</lparam>
<lparam>Address:8855 34901</lparam>
<lparam>Address:8856 34902</lparam>
<lparam>Address:8857 34903</lparam>
<lparam>Address:8858 34904</lparam>
<lparam>Address:8859 34905</lparam>
<lparam>Address:8860 34912</lparam>
<lparam>Address:8861 34913</lparam>
<lparam>Address:8862 34914</lparam>
<lparam>Address:8863 34915</lparam>
<lparam>Address:8864 34916</lparam>
<lparam>Address:8865 34917</lparam>
<lparam>Address:8866 34918</lparam>
<lparam>Address:8867 34919</lparam>
<lparam>Address:8868 34920</lparam>
<lparam>Address:8869 34921</lparam>
<lparam>Address:8870 34928</lparam>
<lparam>Address:8871 34929</lparam>
<lparam>Address:8872 34930</lparam>
<lparam>Address:8873 34931</lparam>
<lparam>Address:8874 34932</lparam>
<lparam>Address:8875 34933</lparam>
<lparam>Address:8876 34934</lparam>
<lparam>Address:8877 34935</lparam>
<lparam>Address:8878 34936</lparam>
<lparam>Address:8879 34937</lparam>
<lparam>Address:8880 34944</lparam>
<lparam>Address:8881 34945</lparam>
<lparam>Address:8882 34946</lparam>
<lparam>Address:8883 34947</lparam>
<lparam>Address:8884 34948</lparam>
<lparam>Address:8885 34949</lparam>
<lparam>Address:8886 34950</lparam>
<lparam>Address:8887 34951</lparam>
<lparam>Address:8888 34952</lparam>
<lparam>Address:8889 34953</lparam>
<lparam>Address:8890 34960</lparam>
<lparam>Address:8891 34961</lparam>
<lparam>Address:8892 34962</lparam>
<lparam>Address:8893 34963</lparam>
<lparam>Address:8894 34964</lparam>
<lparam>Address:8895 34965</lparam>
<lparam>Address:8896 34966</lparam>
<lparam>Address:8897 34967</lparam>
<lparam>Address:8898 34968</lparam>
<lparam>Address:8899 34969</lparam>
<lparam>Address:8900 35072</lparam>
<lparam>Address:8901 35073</lparam>
<lparam>Address:8902 35074</lparam>
<lparam>Address:8903 35075</lparam>
<lparam>Address:8904 35076</lparam>
<lparam>Address:8905 35077</lparam>
<lparam>Address:8906 35078</lparam>
<lparam>Address:8907 35079</lparam>
<lparam>Address:8908 35080</lparam>
<lparam>Address:8909 35081</lparam>
<lparam>Address:8910 35088</lparam>
<lparam>Address:8911 35089</lparam>
<lparam>Address:8912 35090</lparam>
<lparam>Address:8913 35091</lparam>
<lparam>Address:8914 35092</lparam>
<lparam>Address:8915 35093</lparam>
<lparam>Address:8916 35094</lparam>
<lparam>Address:8917 35095</lparam>
<lparam>Address:8918 35096</lparam>
<lparam>Address:8919 35097</lparam>
<lparam>Address:8920 35104</lparam>
<lparam>Address:8921 35105</lparam>
<lparam>Address:8922 35106</lparam>
<lparam>Address:8923 35107</lparam>
<lparam>Address:8924 35108</lparam>
<lparam>Address:8925 35109</lparam>
<lparam>Address:8926 35110</lparam>
<lparam>Address:8927 35111</lparam>
<lparam>Address:8928 35112</lparam>
<lparam>Address:8929 35113</lparam>
<lparam>Address:8930 35120</lparam>
<lparam>Address:8931 35121</lparam>
<lparam>Address:8932 35122</lparam>
<lparam>Address:8933 35123</lparam>
<lparam>Address:8934 35124</lparam>
<lparam>Address:8935 35125</lparam>
<lparam>Address:8936 35126</lparam>
<lparam>Address:8937 35127</lparam>
<lparam>Address:8938 35128</lparam>
<lparam>Address:8939 35129</lparam>
<lparam>Address:8940 35136</lparam>
<lparam>Address:8941 35137</lparam>
<lparam>Address:8942 35138</lparam>
<lparam>Address:8943 35139</lparam>
<lparam>Address:8944 35140</lparam>
<lparam>Address:8945 35141</lparam>
<lparam>Address:8946 35142</lparam>
<lparam>Address:8947 35143</lparam>
<lparam>Address:8948 35144</lparam>
<lparam>Address:8949 35145</lparam>
<lparam>Address:8950 35152</lparam>
<lparam>Address:8951 35153</lparam>
<lparam>Address:8952 35154</lparam>
<lparam>Address:8953 35155</lparam>
<lparam>Address:8954 35156</lparam>
<lparam>Address:8955 35157</lparam>
<lparam>Address:8956 35158</lparam>
<lparam>Address:8957 35159</lparam>
<lparam>Address:8958 35160</lparam>
<lparam>Address:8959 35161</lparam>
<lparam>Address:8960 35168</lparam>
<lparam>Address:8961 35169</lparam>
<lparam>Address:8962 35170</lparam>
<lparam>Address:8963 35171</lparam>
<lparam>Address:8964 35172</lparam>
<lparam>Address:8965 35173</lparam>
<lparam>Address:8966 35174</lparam>
<lparam>Address:8967 35175</lparam>
<lparam>Address:8968 35176</lparam>
<lparam>Address:8969 35177</lparam>
<lparam>Address:8970 35184</lparam>
<lparam>Address:8971 35185</lparam>
<lparam>Address:8972 35186</lparam>
<lparam>Address:8973 35187</lparam>
<lparam>Address:8974 35188</lparam>
<lparam>Address:8975 35189</lparam>
<lparam>Address:8976 35190</lparam>
<lparam>Address:8977 35191</lparam>
<lparam>Address:8978 35192</lparam>
<lparam>Address:8979 35193</lparam>
<lparam>Address:8980 35200</lparam>
<lparam>Address:8981 35201</lparam>
<lparam>Address:8982 35202</lparam>
<lparam>Address:8983 35203</lparam>
<lparam>Address:8984 35204</lparam>
<lparam>Address:8985 35205</lparam>
<lparam>Address:8986 35206</lparam>
<lparam>Address:8987 35207</lparam>
<lparam>Address:8988 35208</lparam>
<lparam>Address:8989 35209</lparam>
<lparam>Address:8990 35216</lparam>
<lparam>Address:8991 35217</lparam>
<lparam>Address:8992 35218</lparam>
<lparam>Address:8993 35219</lparam>
<lparam>Address:8994 35220</lparam>
<lparam>Address:8995 35221</lparam>
<lparam>Address:8996 35222</lparam>
<lparam>Address:8997 35223</lparam>
<lparam>Address:8998 35224</lparam>
<lparam>Address:8999 35225</lparam>
<lparam>Address:9000 32768</lparam></gate>
<gate>
<ID>53</ID>
<type>DE_TO</type>
<position>27,-81</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>54</ID>
<type>BB_CLOCK</type>
<position>50,-90.5</position>
<output>
<ID>CLK</ID>146 </output>
<gparam>angle 180</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>55</ID>
<type>CC_PULSE</type>
<position>-40,-18.5</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AE_OR2</type>
<position>48,-13.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>AE_OR3</type>
<position>17,-40.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>82 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>59</ID>
<type>AM_REGISTER16</type>
<position>-18.5,-92.5</position>
<output>
<ID>OUT_0</ID>115 </output>
<output>
<ID>OUT_1</ID>116 </output>
<output>
<ID>OUT_10</ID>123 </output>
<output>
<ID>OUT_11</ID>124 </output>
<output>
<ID>OUT_12</ID>125 </output>
<output>
<ID>OUT_13</ID>119 </output>
<output>
<ID>OUT_14</ID>120 </output>
<output>
<ID>OUT_15</ID>121 </output>
<output>
<ID>OUT_2</ID>117 </output>
<output>
<ID>OUT_3</ID>113 </output>
<output>
<ID>OUT_4</ID>112 </output>
<output>
<ID>OUT_5</ID>114 </output>
<output>
<ID>OUT_6</ID>118 </output>
<output>
<ID>OUT_7</ID>127 </output>
<output>
<ID>OUT_8</ID>126 </output>
<output>
<ID>OUT_9</ID>122 </output>
<input>
<ID>clear</ID>172 </input>
<input>
<ID>clock</ID>171 </input>
<input>
<ID>count_enable</ID>173 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9001</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>62</ID>
<type>DE_TO</type>
<position>-70,-105</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_AND2</type>
<position>37,-91.5</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_OR2</type>
<position>-84,-105</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>EE_VDD</type>
<position>-18.5,-79</position>
<output>
<ID>OUT_0</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>71</ID>
<type>Pauseulator</type>
<position>-11.5,-108</position>
<input>
<ID>signal</ID>142 </input>
<gparam>angle 0.0</gparam>
<lparam>PAUSE_SIM TRUE</lparam></gate>
<gate>
<ID>77</ID>
<type>CC_PULSE</type>
<position>-41.5,-111.5</position>
<output>
<ID>OUT_0</ID>172 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>GA_LED</type>
<position>-46,-148.5</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AE_OR2</type>
<position>-29,-104</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>CC_PULSE</type>
<position>42,-110.5</position>
<output>
<ID>OUT_0</ID>140 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>84</ID>
<type>BE_JKFF_LOW</type>
<position>44,-101</position>
<input>
<ID>J</ID>140 </input>
<input>
<ID>K</ID>140 </input>
<output>
<ID>Q</ID>139 </output>
<input>
<ID>clock</ID>140 </input>
<output>
<ID>nQ</ID>147 </output>
<gparam>angle 90</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_REGISTER4</type>
<position>-9,-157</position>
<output>
<ID>OUT_0</ID>179 </output>
<output>
<ID>OUT_1</ID>180 </output>
<output>
<ID>OUT_2</ID>181 </output>
<output>
<ID>OUT_3</ID>182 </output>
<input>
<ID>clear</ID>172 </input>
<input>
<ID>clock</ID>195 </input>
<input>
<ID>count_enable</ID>195 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 9</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_REGISTER4</type>
<position>-9,-144</position>
<output>
<ID>OUT_0</ID>183 </output>
<output>
<ID>OUT_1</ID>184 </output>
<output>
<ID>OUT_2</ID>185 </output>
<output>
<ID>OUT_3</ID>186 </output>
<input>
<ID>clear</ID>172 </input>
<input>
<ID>clock</ID>95 </input>
<input>
<ID>count_enable</ID>95 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 9</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_REGISTER4</type>
<position>-8.5,-131.5</position>
<output>
<ID>OUT_0</ID>187 </output>
<output>
<ID>OUT_1</ID>188 </output>
<output>
<ID>OUT_2</ID>189 </output>
<output>
<ID>OUT_3</ID>190 </output>
<input>
<ID>clear</ID>172 </input>
<input>
<ID>clock</ID>197 </input>
<input>
<ID>count_enable</ID>197 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 9</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_REGISTER4</type>
<position>-8.5,-118</position>
<output>
<ID>OUT_0</ID>194 </output>
<output>
<ID>OUT_1</ID>193 </output>
<output>
<ID>OUT_2</ID>192 </output>
<output>
<ID>OUT_3</ID>191 </output>
<output>
<ID>carry_out</ID>142 </output>
<input>
<ID>clear</ID>172 </input>
<input>
<ID>clock</ID>198 </input>
<input>
<ID>count_enable</ID>198 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 9</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_OR2</type>
<position>-22,-164.5</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>195 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AE_OR2</type>
<position>-17.5,-148</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>207 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_OR2</type>
<position>-18,-135.5</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>213 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_OR2</type>
<position>-19,-122</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>210 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>GA_LED</type>
<position>46,-97</position>
<input>
<ID>N_in2</ID>147 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>DE_TO</type>
<position>-77.5,-113.5</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 4</lparam></gate>
<gate>
<ID>101</ID>
<type>AE_SMALL_INVERTER</type>
<position>-85.5,-113.5</position>
<input>
<ID>IN_0</ID>151 </input>
<output>
<ID>OUT_0</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_SMALL_INVERTER</type>
<position>-89.5,-113.5</position>
<input>
<ID>IN_0</ID>150 </input>
<output>
<ID>OUT_0</ID>151 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>103</ID>
<type>AE_SMALL_INVERTER</type>
<position>-93.5,-113.5</position>
<input>
<ID>IN_0</ID>154 </input>
<output>
<ID>OUT_0</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>104</ID>
<type>AE_SMALL_INVERTER</type>
<position>-97.5,-113.5</position>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AE_SMALL_INVERTER</type>
<position>-101.5,-113.5</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>143</ID>
<type>BM_NORX4</type>
<position>15,-155</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>181 </input>
<input>
<ID>IN_2</ID>180 </input>
<input>
<ID>IN_3</ID>179 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>144</ID>
<type>BM_NORX4</type>
<position>15,-142</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>185 </input>
<input>
<ID>IN_2</ID>184 </input>
<input>
<ID>IN_3</ID>183 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>145</ID>
<type>BM_NORX4</type>
<position>15.5,-129.5</position>
<input>
<ID>IN_0</ID>190 </input>
<input>
<ID>IN_1</ID>189 </input>
<input>
<ID>IN_2</ID>188 </input>
<input>
<ID>IN_3</ID>187 </input>
<output>
<ID>OUT</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_REGISTER4</type>
<position>-101,-86.5</position>
<output>
<ID>OUT_0</ID>307 </output>
<input>
<ID>clock</ID>305 </input>
<input>
<ID>count_enable</ID>305 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-118,-2,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_13</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_13</name></connection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-118,-2,-118</points>
<connection>
<GID>90</GID>
<name>OUT_1</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-119,-1,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_12</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_12</name></connection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-119,-1,-119</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-21.5,13,-21.5</points>
<connection>
<GID>1</GID>
<name>OUT_10</name></connection>
<connection>
<GID>12</GID>
<name>IN_10</name></connection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,-162,-10,-162</points>
<intersection>-19 26</intersection>
<intersection>-14 3</intersection>
<intersection>-10 23</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-14,-162,-14,-151.5</points>
<intersection>-162 1</intersection>
<intersection>-151.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-14,-151.5,-9,-151.5</points>
<intersection>-14 3</intersection>
<intersection>-9 24</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-10,-162,-10,-161</points>
<connection>
<GID>87</GID>
<name>clock</name></connection>
<intersection>-162 1</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>-9,-152,-9,-151.5</points>
<connection>
<GID>87</GID>
<name>count_enable</name></connection>
<intersection>-151.5 4</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-19,-164.5,-19,-162</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>-162 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-25.5,13,-25.5</points>
<connection>
<GID>1</GID>
<name>OUT_6</name></connection>
<connection>
<GID>12</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-16.5,13,-16.5</points>
<connection>
<GID>1</GID>
<name>OUT_15</name></connection>
<connection>
<GID>12</GID>
<name>IN_15</name></connection></vsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-15,-135.5,-9.5,-135.5</points>
<connection>
<GID>89</GID>
<name>clock</name></connection>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>-15 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-15,-135.5,-15,-126.5</points>
<intersection>-135.5 1</intersection>
<intersection>-126.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-15,-126.5,-8.5,-126.5</points>
<connection>
<GID>89</GID>
<name>count_enable</name></connection>
<intersection>-15 6</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-42,66.5,-42</points>
<connection>
<GID>23</GID>
<name>carry_in</name></connection>
<connection>
<GID>24</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-122,-16,-112</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>-122 14</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-16,-112,-8.5,-112</points>
<intersection>-16 0</intersection>
<intersection>-8.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-8.5,-113,-8.5,-112</points>
<connection>
<GID>90</GID>
<name>count_enable</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-16,-122,-9.5,-122</points>
<connection>
<GID>90</GID>
<name>clock</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-42,82.5,-42</points>
<connection>
<GID>24</GID>
<name>carry_in</name></connection>
<connection>
<GID>25</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-42,98.5,-42</points>
<connection>
<GID>25</GID>
<name>carry_in</name></connection>
<connection>
<GID>26</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-28.5,13,-28.5</points>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<connection>
<GID>12</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-26.5,13,-26.5</points>
<connection>
<GID>1</GID>
<name>OUT_5</name></connection>
<connection>
<GID>12</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-22.5,13,-22.5</points>
<connection>
<GID>1</GID>
<name>OUT_9</name></connection>
<connection>
<GID>12</GID>
<name>IN_9</name></connection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-19.5,13,-19.5</points>
<connection>
<GID>1</GID>
<name>OUT_12</name></connection>
<connection>
<GID>12</GID>
<name>IN_12</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-23.5,13,-23.5</points>
<connection>
<GID>1</GID>
<name>OUT_8</name></connection>
<connection>
<GID>12</GID>
<name>IN_8</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-20.5,13,-20.5</points>
<connection>
<GID>1</GID>
<name>OUT_11</name></connection>
<connection>
<GID>12</GID>
<name>IN_11</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-30.5,13,-30.5</points>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection>
<connection>
<GID>12</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20.5,-149,18,-149</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<intersection>18 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18,-155,18,-149</points>
<connection>
<GID>143</GID>
<name>OUT</name></connection>
<intersection>-149 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-29.5,13,-29.5</points>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<connection>
<GID>12</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-27.5,13,-27.5</points>
<connection>
<GID>1</GID>
<name>OUT_4</name></connection>
<connection>
<GID>12</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-18.5,13,-18.5</points>
<connection>
<GID>1</GID>
<name>OUT_13</name></connection>
<connection>
<GID>12</GID>
<name>IN_13</name></connection></vsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-22,-123,18.5,-123</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>18.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18.5,-129.5,18.5,-123</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>-123 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-17.5,13,-17.5</points>
<connection>
<GID>1</GID>
<name>OUT_14</name></connection>
<connection>
<GID>12</GID>
<name>IN_14</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-31.5,13,-31.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-24.5,13,-24.5</points>
<connection>
<GID>1</GID>
<name>OUT_7</name></connection>
<connection>
<GID>12</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21,-136.5,18,-136.5</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>18 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18,-142,18,-136.5</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>-136.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120,-104,-87,-104</points>
<connection>
<GID>5</GID>
<name>CLK</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-117 10</intersection>
<intersection>-107.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-107.5,-113.5,-107.5,-104</points>
<intersection>-113.5 21</intersection>
<intersection>-106 19</intersection>
<intersection>-104 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-117,-104,-117,-98</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-107.5,-106,-96,-106</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-107.5 9</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-107.5,-113.5,-103.5,-113.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>-107.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-94.5,13.5,-92</points>
<intersection>-94.5 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-92,13.5,-92</points>
<connection>
<GID>52</GID>
<name>write_enable</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-94.5,15.5,-94.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-5,7.5,-5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-1,7.5,-1</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>9</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-39,104.5,-9</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-9,104.5,-9</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-39,103.5,-8</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-8,103.5,-8</points>
<connection>
<GID>27</GID>
<name>OUT_1</name></connection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-39,102.5,-7</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-7,102.5,-7</points>
<connection>
<GID>27</GID>
<name>OUT_2</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-39,101.5,-6</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-6,101.5,-6</points>
<connection>
<GID>27</GID>
<name>OUT_3</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-39,88.5,-5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-5,88.5,-5</points>
<connection>
<GID>27</GID>
<name>OUT_4</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-39,87.5,-4</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-4,87.5,-4</points>
<connection>
<GID>27</GID>
<name>OUT_5</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-39,86.5,-3</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-3,86.5,-3</points>
<connection>
<GID>27</GID>
<name>OUT_6</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-39,85.5,-2</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-2,85.5,-2</points>
<connection>
<GID>27</GID>
<name>OUT_7</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-39,72.5,-1</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-1,72.5,-1</points>
<connection>
<GID>27</GID>
<name>OUT_8</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-39,71.5,0</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,0,71.5,0</points>
<connection>
<GID>27</GID>
<name>OUT_9</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-39,70.5,1</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,1,70.5,1</points>
<connection>
<GID>27</GID>
<name>OUT_10</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-39,69.5,2</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,2,69.5,2</points>
<connection>
<GID>27</GID>
<name>OUT_11</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-39,56.5,3</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,3,56.5,3</points>
<connection>
<GID>27</GID>
<name>OUT_12</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-39,55.5,4</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,4,55.5,4</points>
<connection>
<GID>27</GID>
<name>OUT_13</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-39,54.5,5</points>
<connection>
<GID>23</GID>
<name>IN_2</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,5,54.5,5</points>
<connection>
<GID>27</GID>
<name>OUT_14</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-39,53.5,6</points>
<connection>
<GID>23</GID>
<name>IN_3</name></connection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,6,53.5,6</points>
<connection>
<GID>27</GID>
<name>OUT_15</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,3,7.5,3</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<connection>
<GID>11</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-39,111.5,-31.5</points>
<connection>
<GID>26</GID>
<name>IN_B_0</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-31.5,111.5,-31.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>37 2</intersection>
<intersection>111.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>37,-31.5,37,-9</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>-31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-39,110.5,-30.5</points>
<connection>
<GID>26</GID>
<name>IN_B_1</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-30.5,110.5,-30.5</points>
<connection>
<GID>12</GID>
<name>OUT_1</name></connection>
<intersection>36.5 3</intersection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36.5,-30.5,36.5,-8</points>
<intersection>-30.5 1</intersection>
<intersection>-8 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36.5,-8,37,-8</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>36.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-39,109.5,-29.5</points>
<connection>
<GID>26</GID>
<name>IN_B_2</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-29.5,109.5,-29.5</points>
<connection>
<GID>12</GID>
<name>OUT_2</name></connection>
<intersection>36 2</intersection>
<intersection>109.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>36,-29.5,36,-7</points>
<intersection>-29.5 1</intersection>
<intersection>-7 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>36,-7,37,-7</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>36 2</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-39,108.5,-28.5</points>
<connection>
<GID>26</GID>
<name>IN_B_3</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-28.5,108.5,-28.5</points>
<connection>
<GID>12</GID>
<name>OUT_3</name></connection>
<intersection>35.5 2</intersection>
<intersection>108.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>35.5,-28.5,35.5,-6</points>
<intersection>-28.5 1</intersection>
<intersection>-6 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>35.5,-6,37,-6</points>
<connection>
<GID>27</GID>
<name>IN_3</name></connection>
<intersection>35.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-39,95.5,-27.5</points>
<connection>
<GID>25</GID>
<name>IN_B_0</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-27.5,95.5,-27.5</points>
<connection>
<GID>12</GID>
<name>OUT_4</name></connection>
<intersection>35 2</intersection>
<intersection>95.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>35,-27.5,35,-5</points>
<intersection>-27.5 1</intersection>
<intersection>-5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>35,-5,37,-5</points>
<connection>
<GID>27</GID>
<name>IN_4</name></connection>
<intersection>35 2</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-39,94.5,-26.5</points>
<connection>
<GID>25</GID>
<name>IN_B_1</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-26.5,94.5,-26.5</points>
<connection>
<GID>12</GID>
<name>OUT_5</name></connection>
<intersection>34.5 2</intersection>
<intersection>94.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>34.5,-26.5,34.5,-4</points>
<intersection>-26.5 1</intersection>
<intersection>-4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>34.5,-4,37,-4</points>
<connection>
<GID>27</GID>
<name>IN_5</name></connection>
<intersection>34.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-39,93.5,-25.5</points>
<connection>
<GID>25</GID>
<name>IN_B_2</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-25.5,93.5,-25.5</points>
<connection>
<GID>12</GID>
<name>OUT_6</name></connection>
<intersection>34 2</intersection>
<intersection>93.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>34,-25.5,34,-3</points>
<intersection>-25.5 1</intersection>
<intersection>-3 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>34,-3,37,-3</points>
<connection>
<GID>27</GID>
<name>IN_6</name></connection>
<intersection>34 2</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-39,92.5,-24.5</points>
<connection>
<GID>25</GID>
<name>IN_B_3</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-24.5,92.5,-24.5</points>
<connection>
<GID>12</GID>
<name>OUT_7</name></connection>
<intersection>33.5 2</intersection>
<intersection>92.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>33.5,-24.5,33.5,-2</points>
<intersection>-24.5 1</intersection>
<intersection>-2 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-2,37,-2</points>
<connection>
<GID>27</GID>
<name>IN_7</name></connection>
<intersection>33.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-39,79.5,-23.5</points>
<connection>
<GID>24</GID>
<name>IN_B_0</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-23.5,79.5,-23.5</points>
<connection>
<GID>12</GID>
<name>OUT_8</name></connection>
<intersection>33 2</intersection>
<intersection>79.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>33,-23.5,33,-1</points>
<intersection>-23.5 1</intersection>
<intersection>-1 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>33,-1,37,-1</points>
<connection>
<GID>27</GID>
<name>IN_8</name></connection>
<intersection>33 2</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-39,78.5,-22.5</points>
<connection>
<GID>24</GID>
<name>IN_B_1</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-22.5,78.5,-22.5</points>
<connection>
<GID>12</GID>
<name>OUT_9</name></connection>
<intersection>32.5 2</intersection>
<intersection>78.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>32.5,-22.5,32.5,0</points>
<intersection>-22.5 1</intersection>
<intersection>0 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>32.5,0,37,0</points>
<connection>
<GID>27</GID>
<name>IN_9</name></connection>
<intersection>32.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-39,77.5,-21.5</points>
<connection>
<GID>24</GID>
<name>IN_B_2</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-21.5,77.5,-21.5</points>
<connection>
<GID>12</GID>
<name>OUT_10</name></connection>
<intersection>32 2</intersection>
<intersection>77.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>32,-21.5,32,1</points>
<intersection>-21.5 1</intersection>
<intersection>1 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>32,1,37,1</points>
<connection>
<GID>27</GID>
<name>IN_10</name></connection>
<intersection>32 2</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-39,76.5,-20.5</points>
<connection>
<GID>24</GID>
<name>IN_B_3</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-20.5,76.5,-20.5</points>
<connection>
<GID>12</GID>
<name>OUT_11</name></connection>
<intersection>31.5 2</intersection>
<intersection>76.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>31.5,-20.5,31.5,2</points>
<intersection>-20.5 1</intersection>
<intersection>2 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>31.5,2,37,2</points>
<connection>
<GID>27</GID>
<name>IN_11</name></connection>
<intersection>31.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-39,63.5,-19.5</points>
<connection>
<GID>23</GID>
<name>IN_B_0</name></connection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-19.5,63.5,-19.5</points>
<connection>
<GID>12</GID>
<name>OUT_12</name></connection>
<intersection>31 2</intersection>
<intersection>63.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>31,-19.5,31,3</points>
<intersection>-19.5 1</intersection>
<intersection>3 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>31,3,37,3</points>
<connection>
<GID>27</GID>
<name>IN_12</name></connection>
<intersection>31 2</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-39,62.5,-18.5</points>
<connection>
<GID>23</GID>
<name>IN_B_1</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-18.5,62.5,-18.5</points>
<connection>
<GID>12</GID>
<name>OUT_13</name></connection>
<intersection>30.5 2</intersection>
<intersection>62.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>30.5,-18.5,30.5,4</points>
<intersection>-18.5 1</intersection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>30.5,4,37,4</points>
<connection>
<GID>27</GID>
<name>IN_13</name></connection>
<intersection>30.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-39,61.5,-17.5</points>
<connection>
<GID>23</GID>
<name>IN_B_2</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-17.5,61.5,-17.5</points>
<connection>
<GID>12</GID>
<name>OUT_14</name></connection>
<intersection>30 4</intersection>
<intersection>61.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30,-17.5,30,5</points>
<intersection>-17.5 1</intersection>
<intersection>5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>30,5,37,5</points>
<connection>
<GID>27</GID>
<name>IN_14</name></connection>
<intersection>30 4</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-39,60.5,-16.5</points>
<connection>
<GID>23</GID>
<name>IN_B_3</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-16.5,60.5,-16.5</points>
<connection>
<GID>12</GID>
<name>OUT_15</name></connection>
<intersection>29.5 2</intersection>
<intersection>60.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>29.5,-16.5,29.5,6</points>
<intersection>-16.5 1</intersection>
<intersection>6 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>29.5,6,37,6</points>
<connection>
<GID>27</GID>
<name>IN_15</name></connection>
<intersection>29.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-57,108,-47</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-57,108,-57</points>
<intersection>-2.5 2</intersection>
<intersection>108 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-2.5,-57,-2.5,-31.5</points>
<intersection>-57 1</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2.5,-31.5,3,-31.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>-2.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-56.5,-3.5,-30.5</points>
<intersection>-56.5 2</intersection>
<intersection>-30.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-3.5,-56.5,107,-56.5</points>
<intersection>-3.5 0</intersection>
<intersection>107 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>107,-56.5,107,-47</points>
<connection>
<GID>26</GID>
<name>OUT_1</name></connection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-3.5,-30.5,3,-30.5</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-56,-4.5,-29.5</points>
<intersection>-56 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-29.5,3,-29.5</points>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4.5,-56,106,-56</points>
<intersection>-4.5 0</intersection>
<intersection>106 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>106,-56,106,-47</points>
<connection>
<GID>26</GID>
<name>OUT_2</name></connection>
<intersection>-56 2</intersection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-55.5,105,-47</points>
<connection>
<GID>26</GID>
<name>OUT_3</name></connection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5.5,-55.5,105,-55.5</points>
<intersection>-5.5 2</intersection>
<intersection>105 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-5.5,-55.5,-5.5,-28.5</points>
<intersection>-55.5 1</intersection>
<intersection>-28.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-5.5,-28.5,3,-28.5</points>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>-5.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-55,92,-47</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6.5,-55,92,-55</points>
<intersection>-6.5 2</intersection>
<intersection>92 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-6.5,-55,-6.5,-27.5</points>
<intersection>-55 1</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-6.5,-27.5,3,-27.5</points>
<connection>
<GID>1</GID>
<name>IN_4</name></connection>
<intersection>-6.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-54.5,91,-47</points>
<connection>
<GID>25</GID>
<name>OUT_1</name></connection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-54.5,91,-54.5</points>
<intersection>-7.5 2</intersection>
<intersection>91 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-7.5,-54.5,-7.5,-26.5</points>
<intersection>-54.5 1</intersection>
<intersection>-26.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-7.5,-26.5,3,-26.5</points>
<connection>
<GID>1</GID>
<name>IN_5</name></connection>
<intersection>-7.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-54,90,-47</points>
<connection>
<GID>25</GID>
<name>OUT_2</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-54,90,-54</points>
<intersection>-8.5 2</intersection>
<intersection>90 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-8.5,-54,-8.5,-25.5</points>
<intersection>-54 1</intersection>
<intersection>-25.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-8.5,-25.5,3,-25.5</points>
<connection>
<GID>1</GID>
<name>IN_6</name></connection>
<intersection>-8.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-53.5,-9.5,-24.5</points>
<intersection>-53.5 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-24.5,3,-24.5</points>
<connection>
<GID>1</GID>
<name>IN_7</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-9.5,-53.5,89,-53.5</points>
<intersection>-9.5 0</intersection>
<intersection>89 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89,-53.5,89,-47</points>
<connection>
<GID>25</GID>
<name>OUT_3</name></connection>
<intersection>-53.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-53,76,-47</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10.5,-53,76,-53</points>
<intersection>-10.5 2</intersection>
<intersection>76 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-10.5,-53,-10.5,-23.5</points>
<intersection>-53 1</intersection>
<intersection>-23.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-10.5,-23.5,3,-23.5</points>
<connection>
<GID>1</GID>
<name>IN_8</name></connection>
<intersection>-10.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-52.5,75,-47</points>
<connection>
<GID>24</GID>
<name>OUT_1</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11.5,-52.5,75,-52.5</points>
<intersection>-11.5 2</intersection>
<intersection>75 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-11.5,-52.5,-11.5,-22.5</points>
<intersection>-52.5 1</intersection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-11.5,-22.5,3,-22.5</points>
<connection>
<GID>1</GID>
<name>IN_9</name></connection>
<intersection>-11.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-52,-12.5,-21.5</points>
<intersection>-52 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,-21.5,3,-21.5</points>
<connection>
<GID>1</GID>
<name>IN_10</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,-52,74,-52</points>
<intersection>-12.5 0</intersection>
<intersection>74 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74,-52,74,-47</points>
<connection>
<GID>24</GID>
<name>OUT_2</name></connection>
<intersection>-52 2</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-51.5,-13.5,-20.5</points>
<intersection>-51.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,-20.5,3,-20.5</points>
<connection>
<GID>1</GID>
<name>IN_11</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,-51.5,73,-51.5</points>
<intersection>-13.5 0</intersection>
<intersection>73 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>73,-51.5,73,-47</points>
<connection>
<GID>24</GID>
<name>OUT_3</name></connection>
<intersection>-51.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-51,-14.5,-19.5</points>
<intersection>-51 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-19.5,3,-19.5</points>
<connection>
<GID>1</GID>
<name>IN_12</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-14.5,-51,60,-51</points>
<intersection>-14.5 0</intersection>
<intersection>60 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60,-51,60,-47</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>-51 2</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-50.5,-15.5,-18.5</points>
<intersection>-50.5 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,-18.5,3,-18.5</points>
<connection>
<GID>1</GID>
<name>IN_13</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15.5,-50.5,59,-50.5</points>
<intersection>-15.5 0</intersection>
<intersection>59 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>59,-50.5,59,-47</points>
<connection>
<GID>23</GID>
<name>OUT_1</name></connection>
<intersection>-50.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-50,-16.5,-17.5</points>
<intersection>-50 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16.5,-17.5,3,-17.5</points>
<connection>
<GID>1</GID>
<name>IN_14</name></connection>
<intersection>-16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-16.5,-50,58,-50</points>
<intersection>-16.5 0</intersection>
<intersection>58 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58,-50,58,-47</points>
<connection>
<GID>23</GID>
<name>OUT_2</name></connection>
<intersection>-50 2</intersection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17.5,-49.5,-17.5,-16.5</points>
<intersection>-49.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17.5,-16.5,3,-16.5</points>
<connection>
<GID>1</GID>
<name>IN_15</name></connection>
<intersection>-17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-17.5,-49.5,57,-49.5</points>
<intersection>-17.5 0</intersection>
<intersection>57 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>57,-49.5,57,-47</points>
<connection>
<GID>23</GID>
<name>OUT_3</name></connection>
<intersection>-49.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-33.5,7,-33.5</points>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<connection>
<GID>13</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-2,-19.5,4</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,4,-18.5,4</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-8.5,-2.5,-7.5</points>
<connection>
<GID>31</GID>
<name>clock</name></connection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-8.5,-2.5,-8.5</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>-2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18.5,6,-18.5,6</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<connection>
<GID>39</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23.5,6,-20.5,6</points>
<connection>
<GID>39</GID>
<name>N_in0</name></connection>
<connection>
<GID>10</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-47,11.5,-33.5</points>
<intersection>-47 5</intersection>
<intersection>-39.5 3</intersection>
<intersection>-33.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>8,-39.5,11.5,-39.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>9,-33.5,11.5,-33.5</points>
<connection>
<GID>1</GID>
<name>clear</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>11.5,-47,23.5,-47</points>
<intersection>11.5 0</intersection>
<intersection>19 29</intersection>
<intersection>23.5 12</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-37.5,-11,51,-11</points>
<connection>
<GID>27</GID>
<name>clear</name></connection>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>-34 9</intersection>
<intersection>-11 15</intersection>
<intersection>-0.5 14</intersection>
<intersection>51 30</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-34,-36,-34,-11</points>
<intersection>-36 11</intersection>
<intersection>-11 7</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-34,-36,23.5,-36</points>
<intersection>-34 9</intersection>
<intersection>23.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>23.5,-47,23.5,-33.5</points>
<intersection>-47 5</intersection>
<intersection>-36 11</intersection>
<intersection>-33.5 28</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-0.5,-11,-0.5,-7.5</points>
<connection>
<GID>31</GID>
<name>clear</name></connection>
<intersection>-11 7</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-11,-11,-11,-9.5</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>-11 7</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>19,-33.5,23.5,-33.5</points>
<connection>
<GID>12</GID>
<name>clear</name></connection>
<intersection>23.5 12</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>19,-47,19,-43.5</points>
<connection>
<GID>58</GID>
<name>IN_2</name></connection>
<intersection>-47 5</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>51,-12.5,51,-11</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>-11 7</intersection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,5,10.5,5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<connection>
<GID>44</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-3,10.5,-3</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-7.5,-11,-7.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,1,10.5,1</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,3.5,-1.5,3.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,5,-12.5,5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<connection>
<GID>35</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>6,-43.5,6,-39.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-92,-106,-92,-106</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,-14.5,7.5,-14.5</points>
<connection>
<GID>1</GID>
<name>load</name></connection>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>7.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>7.5,-14.5,7.5,-9</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14.5,-148,-10,-148</points>
<connection>
<GID>88</GID>
<name>clock</name></connection>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>-14.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-14.5,-148,-14.5,-138.5</points>
<intersection>-148 1</intersection>
<intersection>-138.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-14.5,-138.5,-9,-138.5</points>
<intersection>-14.5 9</intersection>
<intersection>-9 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-9,-139,-9,-138.5</points>
<connection>
<GID>88</GID>
<name>count_enable</name></connection>
<intersection>-138.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,7,7.5,9</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>9 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7.5,9,10.5,9</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-14.5,52,9</points>
<intersection>-14.5 5</intersection>
<intersection>9 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>12.5,-7,12.5,9</points>
<intersection>-7 3</intersection>
<intersection>9 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12.5,9,52,9</points>
<intersection>12.5 1</intersection>
<intersection>22.5 4</intersection>
<intersection>41 7</intersection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>10.5,-7,12.5,-7</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>12.5 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>22.5,7.5,22.5,9</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>9 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>51,-14.5,52,-14.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>41,8,41,9</points>
<connection>
<GID>27</GID>
<name>load</name></connection>
<intersection>9 2</intersection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-46,-36,-13.5</points>
<intersection>-46 3</intersection>
<intersection>-18.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38,-18.5,-36,-18.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-36,-13.5,18,-13.5</points>
<intersection>-36 0</intersection>
<intersection>18 9</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-36,-46,17,-46</points>
<intersection>-36 0</intersection>
<intersection>17 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>17,-46,17,-43.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>-46 3</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>18,-14.5,18,-13.5</points>
<connection>
<GID>12</GID>
<name>count_enable</name></connection>
<intersection>-13.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-6.5,19.5,-6.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-13.5,41,-11</points>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-13.5,45,-13.5</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-37.5,17,-33.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<connection>
<GID>12</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-2.5,19.5,-2.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,1.5,19.5,1.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,3.5,22.5,3.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-4.5,22.5,-4.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-0.5,22.5,-0.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>22.5,-10.5,22.5,-8.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-10.5,22.5,-10.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>22.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-43.5,14.5,5.5</points>
<intersection>-43.5 4</intersection>
<intersection>-14.5 5</intersection>
<intersection>5.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>14.5,5.5,19.5,5.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>14.5,-43.5,15,-43.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>14.5,-14.5,17,-14.5</points>
<connection>
<GID>12</GID>
<name>load</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,-78.5,-100,-78.5</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<connection>
<GID>197</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-96,-5.5,-96</points>
<connection>
<GID>59</GID>
<name>OUT_4</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-90.5,-110,-78.5</points>
<connection>
<GID>201</GID>
<name>CLK</name></connection>
<intersection>-90.5 3</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-110,-78.5,-104,-78.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection>
<intersection>-108 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110,-90.5,-102,-90.5</points>
<connection>
<GID>191</GID>
<name>clock</name></connection>
<intersection>-110 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-108,-81.5,-108,-78.5</points>
<intersection>-81.5 5</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-108,-81.5,-101,-81.5</points>
<connection>
<GID>191</GID>
<name>count_enable</name></connection>
<intersection>-108 4</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-97,-5.5,-97</points>
<connection>
<GID>59</GID>
<name>OUT_3</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-95,-5.5,-95</points>
<connection>
<GID>59</GID>
<name>OUT_5</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-87.5,-92.5,-87.5</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<connection>
<GID>207</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-100,-5.5,-100</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-99,-5.5,-99</points>
<connection>
<GID>59</GID>
<name>OUT_1</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96,-78.5,-96,-78.5</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<connection>
<GID>208</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-98,-5.5,-98</points>
<connection>
<GID>59</GID>
<name>OUT_2</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-94,-5.5,-94</points>
<connection>
<GID>59</GID>
<name>OUT_6</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-87,-5.5,-87</points>
<connection>
<GID>59</GID>
<name>OUT_13</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_13</name></connection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-86,-5.5,-86</points>
<connection>
<GID>59</GID>
<name>OUT_14</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_14</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-85,-5.5,-85</points>
<connection>
<GID>59</GID>
<name>OUT_15</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_15</name></connection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-92,-78.5,-92,-78.5</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<connection>
<GID>212</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-91,-5.5,-91</points>
<connection>
<GID>59</GID>
<name>OUT_9</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_9</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-90,-5.5,-90</points>
<connection>
<GID>59</GID>
<name>OUT_10</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_10</name></connection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88,-78.5,-88,-78.5</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<connection>
<GID>213</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-89,-5.5,-89</points>
<connection>
<GID>59</GID>
<name>OUT_11</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_11</name></connection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84,-78.5,-84,-78.5</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<connection>
<GID>215</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-88,-5.5,-88</points>
<connection>
<GID>59</GID>
<name>OUT_12</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_12</name></connection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80,-78.5,-66,-78.5</points>
<connection>
<GID>215</GID>
<name>OUT_0</name></connection>
<connection>
<GID>206</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-92,-5.5,-92</points>
<connection>
<GID>59</GID>
<name>OUT_8</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_8</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-93,-5.5,-93</points>
<connection>
<GID>59</GID>
<name>OUT_7</name></connection>
<connection>
<GID>52</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88,-106,-87,-106</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-34.5,-173,33,-173</points>
<intersection>-34.5 11</intersection>
<intersection>-25 25</intersection>
<intersection>33 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>33,-173,33,-91</points>
<intersection>-173 5</intersection>
<intersection>-91.5 14</intersection>
<intersection>-91 46</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-34.5,-173,-34.5,-103</points>
<intersection>-173 5</intersection>
<intersection>-103 24</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>33,-91.5,34,-91.5</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<intersection>33 6</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-34.5,-103,-32,-103</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>-34.5 11</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>-25,-173,-25,-165.5</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>-173 5</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>12.5,-91,33,-91</points>
<connection>
<GID>52</GID>
<name>write_clock</name></connection>
<intersection>27 50</intersection>
<intersection>33 6</intersection></hsegment>
<vsegment>
<ID>50</ID>
<points>27,-91,27,-83</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-91 46</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-81,-105,-72,-105</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<connection>
<GID>62</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-98,42,-92.5</points>
<connection>
<GID>84</GID>
<name>Q</name></connection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-92.5,42,-92.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>42,-104,46,-104</points>
<connection>
<GID>84</GID>
<name>K</name></connection>
<connection>
<GID>84</GID>
<name>clock</name></connection>
<connection>
<GID>84</GID>
<name>J</name></connection>
<intersection>42 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>42,-108.5,42,-104</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>-104 3</intersection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,-113,-6.5,-108</points>
<connection>
<GID>71</GID>
<name>signal</name></connection>
<connection>
<GID>90</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-90.5,46,-90.5</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<connection>
<GID>54</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-98,46,-98</points>
<connection>
<GID>84</GID>
<name>nQ</name></connection>
<connection>
<GID>96</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-91.5,-113.5,-91.5,-113.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-113.5,-87.5,-113.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-83.5,-113.5,-79.5,-113.5</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<connection>
<GID>97</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-99.5,-113.5,-99.5,-113.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-95.5,-113.5,-95.5,-113.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-104,-19.5,-102</points>
<connection>
<GID>59</GID>
<name>clock</name></connection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26,-104,-19.5,-104</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>-19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39.5,-111.5,-17.5,-111.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>-32 16</intersection>
<intersection>-17.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-17.5,-111.5,-17.5,-102</points>
<connection>
<GID>59</GID>
<name>clear</name></connection>
<intersection>-111.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-32,-171,-32,-105</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>-171 23</intersection>
<intersection>-163.5 26</intersection>
<intersection>-147 38</intersection>
<intersection>-134.5 18</intersection>
<intersection>-121 19</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-32,-134.5,-21,-134.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>-32 16</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-32,-121,-22,-121</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-32 16</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-32,-171,-1.5,-171</points>
<intersection>-32 16</intersection>
<intersection>-1.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>-1.5,-171,-1.5,-122</points>
<intersection>-171 23</intersection>
<intersection>-161 37</intersection>
<intersection>-148 34</intersection>
<intersection>-135.5 35</intersection>
<intersection>-122 36</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>-32,-163.5,-25,-163.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-32 16</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>-8,-148,-1.5,-148</points>
<connection>
<GID>88</GID>
<name>clear</name></connection>
<intersection>-1.5 24</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>-7.5,-135.5,-1.5,-135.5</points>
<connection>
<GID>89</GID>
<name>clear</name></connection>
<intersection>-1.5 24</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>-7.5,-122,-1.5,-122</points>
<connection>
<GID>90</GID>
<name>clear</name></connection>
<intersection>-1.5 24</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-8,-161,-1.5,-161</points>
<connection>
<GID>87</GID>
<name>clear</name></connection>
<intersection>-1.5 24</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>-32,-147,-20.5,-147</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>-32 16</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18.5,-83,-18.5,-80</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<connection>
<GID>59</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-158,11,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_0</name></connection>
<intersection>-158 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-158,12,-158</points>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<connection>
<GID>143</GID>
<name>IN_3</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-157,10,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_1</name></connection>
<intersection>-157 1</intersection>
<intersection>-156 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-157,10,-157</points>
<connection>
<GID>87</GID>
<name>OUT_1</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>10,-156,12,-156</points>
<connection>
<GID>143</GID>
<name>IN_2</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-156,9,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_2</name></connection>
<intersection>-156 1</intersection>
<intersection>-154 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-156,9,-156</points>
<connection>
<GID>87</GID>
<name>OUT_2</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>9,-154,12,-154</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-155,8,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_3</name></connection>
<intersection>-155 1</intersection>
<intersection>-152 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-155,8,-155</points>
<connection>
<GID>87</GID>
<name>OUT_3</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>8,-152,12,-152</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-145,7,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_4</name></connection>
<intersection>-145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-145,12,-145</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<connection>
<GID>144</GID>
<name>IN_3</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-5,-144,6,-144</points>
<connection>
<GID>88</GID>
<name>OUT_1</name></connection>
<intersection>6 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>6,-144,6,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_5</name></connection>
<intersection>-144 3</intersection>
<intersection>-143 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6,-143,12,-143</points>
<connection>
<GID>144</GID>
<name>IN_2</name></connection>
<intersection>6 4</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5,-143,5,-143</points>
<connection>
<GID>88</GID>
<name>OUT_2</name></connection>
<intersection>5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>5,-143,5,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_6</name></connection>
<intersection>-143 1</intersection>
<intersection>-141 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>5,-141,12,-141</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>5 3</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-5,-142,4,-142</points>
<connection>
<GID>88</GID>
<name>OUT_3</name></connection>
<intersection>4 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>4,-142,4,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_7</name></connection>
<intersection>-142 3</intersection>
<intersection>-139 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>4,-139,12,-139</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>4 4</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-132.5,3,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_8</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_8</name></connection>
<intersection>-132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-132.5,12.5,-132.5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<connection>
<GID>145</GID>
<name>IN_3</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-131.5,2,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_9</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_9</name></connection>
<intersection>-131.5 1</intersection>
<intersection>-130.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-131.5,2,-131.5</points>
<connection>
<GID>89</GID>
<name>OUT_1</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2,-130.5,12.5,-130.5</points>
<connection>
<GID>145</GID>
<name>IN_2</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-130.5,1,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_10</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_10</name></connection>
<intersection>-130.5 1</intersection>
<intersection>-128.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-130.5,1,-130.5</points>
<connection>
<GID>89</GID>
<name>OUT_2</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,-128.5,12.5,-128.5</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-129.5,0,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_11</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_11</name></connection>
<intersection>-129.5 1</intersection>
<intersection>-126.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-129.5,0,-129.5</points>
<connection>
<GID>89</GID>
<name>OUT_3</name></connection>
<intersection>0 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,-126.5,12.5,-126.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-116,-4,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_15</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_15</name></connection>
<intersection>-116 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-116,-4,-116</points>
<connection>
<GID>90</GID>
<name>OUT_3</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-117,-3,-103.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_14</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_14</name></connection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-117,-3,-117</points>
<connection>
<GID>90</GID>
<name>OUT_2</name></connection>
<intersection>-3 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 1>
<page 2>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 2>
<page 3>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 3>
<page 4>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 4>
<page 5>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 5>
<page 6>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 6>
<page 7>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 7>
<page 8>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 8>
<page 9>
<PageViewport>0,384.093,1224,-220.907</PageViewport></page 9></circuit>